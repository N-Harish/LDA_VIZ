��V�      ]�(]�(K K��KK��KK��KK��KK��KK��KK��KK��KK��K	K��K
K��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��K K��K!K��K"K��K#K��K$K��K%K��K&K��K'K��K(K��K)K��K*K��K+K��K,K��K-K��K.K��K/K��K0K��K1K��K2K��K3K��K4K��K5K��K6K��K7K��K8K��K9K��K:K��K;K��K<K��K=K��K>K��K?K��K@K��KAK��KBK��KCK��KDK��KEK��KFK��KGK��KHK��KIK��KJK��KKK��KLK��KMK��KNK��KOK��KPK��KQK��KRK��KSK��KTK��KUK��KVK��KWK��KXK��KYK��KZK��K[K��K\K��K]K��K^K��K_K��K`K��KaK��KbK��KcK��KdK��KeK��KfK��KgK��KhK��KiK��KjK��KkK	��KlK��KmK��KnK��KoK��KpK��KqK��KrK��KsK��KtK��KuK��KvK��KwK��KxK��KyK��KzK��K{K��K|K��K}K��K~K��KK��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K
��K�K��K�K��K�K��K�K��K�K��K�K	��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K	��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK"��MJK	��MKK��MLK��MMK	��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K
��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK
��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K"��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK&��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK
��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K(��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK
��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK%��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK	��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K#��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��e(M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K
��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K
��M9K��M:K��M;K��M<K��M=K��M>K
��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK
��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK9��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K"��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK
��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK	��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K
��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K&��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK
��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K	��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK
��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK	��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��e(M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK	��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK	��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK	��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��e]�(KK��KK��KK��KK	��KK��K	K��K
K��KK��KK��KK��KK��KK��KK��KK��KK��K!K��K$K��K%K��K)K��K*K��K,K��K-K��K.K��K0K��K3K��K4K��K8K��K9K��K:K��K=K��K?K��K@K��KAK��KCK��KDK��KEK��KFK��KHK��KJK��KLK��KOK��KPK��KRK��KSK��KTK
��KUK��KVK��KXK��KYK��KZK��K[K��K\K��K^K��K`K��KcK��KdK��KgK��KkK��KlK��KnK��KrK��KtK��KvK��KwK��KxK��K{K��K|K��K�K!��K�K��K�K��K�K��K�K��K�K��K�K	��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M"K��M&K��M'K��M,K��M-K��M.K��M1K��M2K��M3K��M5K&��M7K��M;K��M=K	��M>K
��MDK��MFK��MHK��MIK��MJK	��MKK��MLK��MMK��MOK��MUK��MVK��MWK��MYK��MZK	��M[K��M\K��MaK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MmK��MnK��MpK��MqK��MrK��MuK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M K��M
K��MK��MK	��MK��MK��MK��MK��MK��MK��MK��MK��M K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M+K��M,K��M.K��M/K��M4K��M6K��M<K��M=K��M@K��MAK��MDK��MHK��MMK��MPK��MQK��MRK��MUK��MXK��M\K��M]K��MbK��McK��MdK��MfK��MgK��MhK��MiK��MjK��MnK��MpK��MrK��MwK��MxK��MyK��MzK��M{K��M|K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK
��M!K��M#K��M$K��M%K��M&K��M'K��M(K��M*K��M.K��M0K��M1K��M3K��M4K��M6K��M7K��M8K��M<K��MBK��MCK��MDK��MHK��MJK��MKK��MNK��MSK��MYK��MZK��M\K��M]K��M_K��MbK	��McK��MdK��MeK��MfK��MgK��MjK��MnK��MrK��MuK��MvK��MwK��M{K��M~K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K	��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M"K��M#K��M)K��M,K��M1K��M4K��M5K��M6K��M8K��M9K��M<K��M=K��M>K��M?K��M@K��MBK��MCK��MDK��MEK��MGK��MJK��MLK��MMK��MNK
��MQK��MRK��MUK��MVK��MXK��MYK��MZK��M\K��M_K��MaK��MbK	��McK��MfK��MgK��MiK%��MjK��MuK��MwK��MxK��MyK��MzK��M}K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K*��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��MK
��MK��MK��MK��M	K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M$K��M'K��M(K��M*K��M+K��M-K��M0K��M1K��M2K��M3K��M5K��M7K��M8K��M;K��M>K��M?K��M@K��MAK��MDK��MEK��MFK��MNK��MPK��MQK��MUK	��MWK��MYK��MZK��M\K
��M]K��M_K��M`K��MaK��MeK��MfK��MkK��MmK��MrK��MsK��MtK��MuK��MwK��MzK��M}K��MK��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K	��MK��MK
��MK	��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK	��MK��MK��MK��MK��M K��M!K��M%K��M(K��M)K��M*K��M+K	��M-K��M.K��M0K��M1K��M2K��M5K��M7K��M8K��M;K��M<K��M>K��M@K��MAK��MCK��MEK��MFK��MGK��MHK��MLK��MNK
��MQK
��MRK��MSK��MWK��MXK��MZK��M]K��M^K��M_K��M`K��MbK��McK��MdK��MeK��MhK
��MjK��MkK��MlK��MoK��MpK��MqK
��MwK��MzK��M{K��M|K��M}K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M#K��M$K��M%K��M&K��M'K��M(K��M/K��M0K��M1K��M5K��M6K��M8K��M:K��M<K��M=K��M?K��MAK��MBK��MCK��MDK��MEK��MHK��MIK��MKK��MNK��MOK��MQK��MRK��MSK��MTK��MUK��MVK��MWK	��MXK��MZK��M\K��M]K��M_K��M`K��MbK��MdK��MgK��MiK��MmK��MoK��MpK��MrK��MtK��MuK��MwK��MxK��MyK��M{K��M|K��M~K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��e(M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK
��MK��MK��MK��MK��MK��MK��M K��M"K��M&K��M'K��M(K��M*K��M.K��M/K��M0K��M3K��M5K��M6K��M7K��M8K��M<K,��M?K��M@K��MBK��MFK��MLK��MMK��MNK��MQK��MRK��MTK��MVK��MWK��M\K��M^K��M_K��M`K��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MsK��MvK��MxK��MyK
��MzK��M{K	��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K/��M�K��M�K��M�K��M�K%��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M 	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M		K��M
	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M 	K��M!	K��M"	K��M#	K��M$	K��M%	K��M&	K��M'	K��M(	K��M)	K��M*	K��M+	K��M,	K��M-	K��M.	K��M/	K��M0	K��M1	K��M2	K��M3	K��M4	K��M5	K��M6	K��M7	K��M8	K��M9	K��M:	K��M;	K��M<	K��M=	K��M>	K��M?	K��M@	K��MA	K��MB	K��MC	K��MD	K��ME	K��MF	K��MG	K��MH	K��MI	K��MJ	K��MK	K��ML	K��MM	K��MN	K��MO	K��MP	K��MQ	K��MR	K��MS	K��MT	K��MU	K��MV	K��MW	K��MX	K��MY	K��MZ	K��M[	K��M\	K��M]	K��M^	K��M_	K��M`	K��Ma	K��Mb	K��Mc	K��Md	K��Me	K��Mf	K��Mg	K��Mh	K��Mi	K��Mj	K��Mk	K��Ml	K��Mm	K��Mn	K��Mo	K��Mp	K��Mq	K��Mr	K��Ms	K��Mt	K��Mu	K��Mv	K��Mw	K��Mx	K��My	K��Mz	K��M{	K��M|	K��M}	K��M~	K��M	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M 
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M	
K��M

K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M 
K��M!
K��M"
K��M#
K��M$
K��M%
K��M&
K��M'
K��M(
K��M)
K��M*
K��M+
K��M,
K��M-
K��M.
K��M/
K��M0
K��M1
K��M2
K��M3
K��M4
K��M5
K��M6
K��M7
K��M8
K��M9
K��M:
K��M;
K��M<
K��M=
K��M>
K��M?
K��M@
K��MA
K��MB
K��MC
K��MD
K��ME
K��MF
K��MG
K��MH
K��MI
K��MJ
K��MK
K��ML
K��MM
K��MN
K��MO
K��MP
K��MQ
K��MR
K��MS
K��MT
K��MU
K��MV
K��MW
K��MX
K��MY
K��MZ
K��M[
K��M\
K��M]
K��M^
K��M_
K��M`
K��Ma
K��Mb
K��Mc
K��Md
K��Me
K��Mf
K��Mg
K��Mh
K��Mi
K��Mj
K��Mk
K��Ml
K��Mm
K��Mn
K��Mo
K��Mp
K��Mq
K��Mr
K��Ms
K��Mt
K��Mu
K��Mv
K��Mw
K��Mx
K��My
K��Mz
K��M{
K��M|
K��M}
K��M~
K��M
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��e(MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK	��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��e]�(KK��KK��KK��KK��K	K��K
K��KK��KK��KK��KK
��KK��KK��KK��KK��KK��KK��KK��KK��K!K��K$K��K'K��K)K��K*K��K,K��K-K	��K.K��K3K��K4K��K7K��K8K��K9K��K:K��K=K��K>K��K?K��K@K��KCK��KDK��KEK��KFK��KHK��KIK��KKK��KOK��KPK��KQK��KRK��KTK��KUK��KVK��K[K��K\K��K^K��K_K��K`K��KaK��KbK��KdK��KfK��KjK��KkK	��KlK��KmK��KnK��KqK��KrK��KtK	��KuK��KvK��KwK��KxK��KyK��KzK��K{K��K|K��K}K��K~K��KK��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K
��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K	��K�K	��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K	��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��MK��MK��MK��MK��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK	��MK��M K��M"K��M#K��M&K��M'K��M(K��M*K��M+K��M,K��M-K��M/K��M1K��M2K��M3K��M5K��M6K��M7K��M8K��M;K��M=K��M>K��MAK��MBK��MDK��MEK��MFK��MGK��MHK��MIKB��MJK��MKK��MLK��MMK��MOK��MRK��MUK��MWK��MYK��MZK��M[K��M\K��M]K��MaK��MdK��MhK��MjK��MkK��MmK��MnK��MpK��MqK��MrK��MsK��MuK��MvK��MyK��MzK��M{K��M|K��M}K��MK��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K%��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K!��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��MK��M	K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M"K��M$K��M%K��M&K��M'K	��M(K��M+K��M,K��M.K��M4K��M6K��M8K��M<K��M@K��MAK��MDK��MFK��MHK��MIK��MJK��MLK��MMK��MPK��MQK��MRK��MSK��MXK��MYK��M\K��M]K��M_K��M`K��MbK��McK��MdK��MfK��MgK��MiK��MnK��MrK��MsK��MxK��MyK��M{K��M|K��M~K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M!K��M#K��M$K��M'K��M,K��M.K��M0K��M2K��M3K��M4K��M6K��M:K��M<K��M=K��M?K��MBK��MCK��MDK��MFK��MHK��MJK��MKK��MNK��MSK��MTK��MVK��MXK��MYK��MZK��M\K��M_K��MaK��MbK��McK��MfK��MgK��MiK��MjK��MnK��MoK��MrK��MuK��MwK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��M K��M"K��M#K��M%K��M)K��M,K��M1K��M5K��M6K��M7K��M8K��M9K��M:K��M<K��M=K��M>K��M?K��MBK��MCK��MDK��MEK	��MGK��MHK��MIK��MJK��MLK��MRK��MSK��MTK��MUK��MVK��MYK��MZK��M[K��M\K��M_K��MaK��MbK��McK	��MdK��MeK��MfK��MhK��MiK��MkK��MnK��MoK��MuK��MvK��MxK��MzK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK
��MK��MK��MK��MK��MK��MK��M K��M!K	��M"K��M#K��M$K��M%K��M'K��M(K��M*K��M+K��M,K��M0K��M1K��M2K��M3K��M5K��M6K��M7K��M8K��M;K��M>K��M?K��M@K��MAK��MCK��MDK��MEK��MFK��MIK��MOK��MPK��MQK��MRK��MUK��MWK��MYK��M\K��M_K��M`K��MaK��MbK��MdK��MeK��MfK��MhK��MmK��MpK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MzK��M}K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK
��MK��MK��M K��M!K��M%K��M&K��M(K��M)K��M*K��M+K	��M-K��M/K��M0K��M2K��M5K��M6K��M7K��M8K��M9K��M;K��M<K��M>K��M?K��MAK��MBK��MCK��MEK��MFK��MGK��MLK��MNK��MQK	��MRK��MTK��MUK��MVK��MWK��MZK��M[K��M]K��M^K��M_K��MbK��McK��MdK��MhK��MjK��MlK��MpK��MqK��MtK��MwK��MzK
��M{K��M}K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M#K��M$K��M%K��M&K��M'K��M(K��M+K��M0K��M1K��M6K��M<K��MBK��MDK��MEK��MHK��MIK��MLK��MOK��MQK��MSK��MTK��MUK��MWK��MXK��M\K��M]K��M_K��MaK��MbK��MeK��MfK��MgK��MiK��MoK��MrK��MtK��MvK��e(MwK��MxK��MyK��M{K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M$K��M%K��M&K��M(K��M*K��M.K��M/K��M0K��M3K��M7K��M:K��M<K��M>K��MAK��MBK��MEK��MFK��MGK��MIK��MMK��MQK��MRK��MTK��MVK��MZK��M]K��M^K��M_K��McK��MeK��MfK��MgK��MhK��MjK ��MoK��MtK��MwK��MyK��MzK��M{K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M	K
��M!	K��M#	K��M$	K��M&	K��M*	K��M+	K��M.	K��M8	K��M<	K��MB	K��ME	K��MF	K��MG	K��MJ	K��MK	K��MR	K��MS	K��MT	K��MZ	K��M[	K��M\	K��Ma	K��Mc	K��Md	K��Mf	K��Mg	K��Mi	K��Ml	K��Mn	K��Mr	K��Ms	K��Mu	K��Mv	K��My	K��Mz	K��M|	K��M}	K��M~	K��M	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M
K��M	
K��M
K��M
K��M
K��M
K��M
K��M 
K��M"
K��M#
K��M&
K��M-
K��M.
K��M/
K��M1
K��M5
K��M:
K��M;
K��M<
K��M?
K��MB
K��MI
K��MK
K��ML
K��MM
K��MT
K��MV
K��MY
K��M\
K��M]
K��Mb
K��Ml
K��Mm
K��M|
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M#K��M%K��M&K��M'K��M+K��M/K��M0K��M2K��M3K��M5K��M6K��M8K��MDK��MHK��MIK��MMK��MRK��MVK��MaK��MfK��MgK��MiK��MqK��MrK��MuK��MvK��MwK��MxK��MyK��M{K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M#K��M'K��M*K��M-K��M6K��M7K��M9K��M;K��M=K��M?K��MEK��MMK��MPK��MSK��MTK��MUK��MVK��M[K��M]K��MgK��MhK��MlK��MvK��MzK��M{K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��e(MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��e]�(KK��KK��KK��KK��KK��K	K��K
K��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��KK��K!K��K%K��K(K��K)K��K*K��K-K��K.K��K0K��K1K��K2K��K3K��K4K��K7K��K8K��K9K��K:K��K<K��K=K��K>K��K?K��K@K��KCK��KDK��KEK��KJK��KKK��KOK��KPK��KRK��KTK��KUK��KXK��KYK��KZK��K[K��K\K
��K^K��K`K��KaK��KbK��KcK��KdK��KgK��KhK��KjK��KkK��KlK��KmK��KnK��KsK��KtK��KuK��KvK��KwK��KxK��KyK��KzK��K{K��K|K��K~K��KK��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��K�K��MK��MK	��MK��MK��MK	��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M"K��M&K��M'K��M-K��M.K��M1K��M2K��M3K��M5KN��M7K��M;K��M=K��M>K��MBK��MDK��MEK��MFK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MQK��MRK��MUK��MWK��MYK��MZK��M[K��M\K��MaK��MbK��MdK��MfK��MhK��MjK��MkK��MmK
��MnK��MpK��MrK��MsK��MuK��MvK��MyK��MzK��M|K��M}K��M~K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K!��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K"��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��M K��M"K��M%K��M&K��M'K��M+K��M,K��M.K��M6K��M=K��M@K��MAK��MDK��MFK��MHK��MIK��MJK��MLK��MMK��MOK��MPK	��MQK��MRK��MSK��MXK��M\K��MbK��McK��MdK��MfK��MgK��MiK��MnK��MqK��MrK��MsK��MwK��MxK��M{K��M|K��M~K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M!K��M#K��M$K��M%K��M&K��M'K��M(K��M+K��M.K��M0K��M1K��M3K��M4K��M6K��M<K
��M=K��M@K��MBK��MCK��MFK��MHK��MIK��MJK��MKK��MNK��MSK��MYK��MZK��M_K��MaK��MbK��McK��MfK��MgK��MjK��MlK��MnK��MuK��MvK��MwK��M~K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M"K��M#K��M$K��M%K��M'K��M)K��M,K��M1K��M2K��M5K��M6K��M8K��M9K��M:K��M=K��M>K��M?K��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MNK��MOK��MPK��MUK��MVK��MYK��MZK��M[K��M\K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MiK��MkK��MnK��MqK��MtK��MuK��MwK��MxK��MyK��MzK��M}K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K
��M$K��M'K��M(K��M+K��M,K��M.K��M0K��M1K��M3K��M5K��M6K��M7K��M8K
��M:K��M=K��M>K ��M?K��M@K��MAK��MCK��MDK��MEK��MFK��MJK��MLK��MMK��MNK��MOK��MQK��MUK(��MYK	��M\K��M^K��M_K	��M`K��MaK��MbK��McK��MeK��MfK	��MjK��MkK��MmK��MpK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MzK��M}K��MK��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�Kӆ�M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK*��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M#K��M%K��M&K��M(K��M)K��M*K��M+K��M-K��M/K��M0K��M2K��M5K��M7K��M8K��M;K��M<K��M>K��M@K��MBK��MCK��MDK��MEK��MFK
��MGK��MJK��MLK��MMK��MNK��MPK��MQK��MRK��MVK��MWK��MYK��MZK��M[K��M]K��M^K��M_K��M`K��MbK��McK��MeK��MhK��MjK��MkK��MlK��MpK��MqK	��MuK��MwK��MzK
��M{K��M|K��M}K��M~K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K	��M�K��M�K��M�K��M�K��M�K
��M K��MK��MK��MK��MK��MK��MK	��M	K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M#K��M$K��M%K��M&K��M'K��M(K��M+K��M.K��M0K��M1K��M6K��M<K��MBK��MDK��MFK��MGK��MIK��MOK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M]K��M_K
��M`K��MbK��MdK��MeK��MfK��MgK��MnK��MoK��MpK��MrK��MtK��MwK��MxK��e(MyK	��M{K��M|K��M}K��M~K	��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K
��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M%K��M&K	��M'K��M(K��M,K��M/K��M0K��M2K��M3K��M6K��M7K��M:K��M<K��M@K��MAK��MDK��MFK��MLK��MMK��MPK��MQK��MVK��M[K��M]K��M_K��MeK��MfK��MgK��MhK��MjK&��MkK��MlK��MoK��MrK��MuK��MvK��MyK��MzK��M{K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M	K��M	K��M	K��M	K��M	K��M	K��M	K��M"	K��M$	K��M+	K��M,	K��M9	K��M<	K��M?	K��MF	K��MM	K��MN	K��MR	K��MT	K��MZ	K��M[	K��M`	K��Ma	K��Md	K��Mf	K��Ml	K��Mn	K��My	K��Mz	K��M}	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M�	K��M
K��M	
K��M
K��M
K��M
K��M
K��M
K��M
K��M
K��M 
K��M#
K��M%
K��M&
K��M,
K��M-
K��M.
K��M:
K��M;
K��M?
K��MC
K��ME
K��MG
K��MK
K��MS
K��MV
K��MW
K��MX
K��M\
K��Ml
K��M{
K��M|
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M�
K��M K��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK
��M!K��M#K��M$K��M&K��M)K��M/K��M0K��M5K��M6K��M8K��MBK��MCK��MEK��MFK��MGK��MHK��MIK��MJK��MOK��MPK��MQK��MRK��M^K��MaK��McK��MeK��MgK��MiK��MjK��MnK��MpK��MsK��MuK��MxK��MyK��M{K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��M
K��MK��MK��MK��MK��MK��MK��MK��M!K��M#K��M)K��M*K��M-K��M?K��MEK��MOK��MQK��MTK��MUK��MZK��M[K��M]K��M^K��MbK��MhK��MvK��MwK��MzK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M-K��M4K��M;K��MOK��MRK��MXK��M\K��M`K��McK��MhK��MsK��MvK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��M	K��MK��MK��M*K��MJK��MQK��MSK��MTK��MXK��MZK��M]K��M`K��MlK��MmK��MqK��MrK��M}K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��MK��MK��MK��M K��M&K��M'K��M)K��M2K��M4K��M6K��M7K��M9K��MBK��MKK��MUK��MVK��MWK��M_K��MaK��MiK��MoK��MpK��MrK��MtK��MuK��MwK��MxK��M|K��M}K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��M#K��M$K��M,K��M3K��M6K��M9K��M>K��M?K��MDK��MFK��MHK��MKK��MYK��MfK��MgK��MoK��MsK��MvK��MzK��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��e(M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M K��MK��MK��MK��MK��MK��MK��MK��MK��M	K��M
K��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��MK��M K��M!K��M"K��M#K��M$K��M%K��M&K��M'K��M(K��M)K��M*K��M+K��M,K��M-K��M.K��M/K��M0K��M1K��M2K��M3K��M4K��M5K��M6K��M7K��M8K��M9K��M:K��M;K��M<K��M=K��M>K��M?K��M@K��MAK��MBK��MCK��MDK��MEK��MFK��MGK��MHK��MIK��MJK��MKK��MLK��MMK��MNK��MOK��MPK��MQK��MRK��MSK��MTK��MUK��MVK��MWK��MXK��MYK��MZK��M[K��M\K��M]K��M^K��M_K��M`K��MaK��MbK��McK��MdK��MeK��MfK��MgK��MhK��MiK��MjK��MkK��MlK��MmK��MnK��MoK��MpK��MqK��MrK��MsK��MtK��MuK��MvK��MwK��MxK��MyK��MzK��M{K��M|K��M}K��M~K��MK��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��M�K��ee.