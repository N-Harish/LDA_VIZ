�cgensim.corpora.dictionary
Dictionary
q )�q}q(X   token2idq}q(X   abilityqK X	   abolitionqKX   absentqKX   abuseqKX   acceptq	KX   accessq
KX   accidentqKX
   accidentalqKX   accountqKX   accuseqK	X   actionqK
X   activistqKX   activityqKX   actressqKX   addqKX   addressqKX   adelaideqKX   adjournqKX   administratorqKX   admitqKX   advanceqKX	   advantageqKX	   adventureqKX   adviceqKX   adviseqKX   advocateqKX   affairqKX   affectq KX	   affectingq!KX   affordq"KX
   affordableq#KX   afghanq$KX   afraidq%K X   africanq&K!X   afridiq'K"X   agassisq(K#X   agencyq)K$X   agendaq*K%X   agentq+K&X   agforceq,K'X
   aggressionq-K(X   agreeq.K)X	   agreementq/K*X   agriculturalq0K+X   agricultureq1K,X   aheadq2K-X   aimq3K.X   airq4K/X   aircraftq5K0X   aireq6K1X   airliftq7K2X   airlineq8K3X   airportq9K4X   akbarq:K5X   alainq;K6X   alarmq<K7X   alcoholq=K8X   alertq>K9X   aliceq?K:X   alienateq@K;X   alightqAK<X   aliveqBK=X
   allegationqCK>X   allegeqDK?X   allegedqEK@X   allianceqFKAX   allocateqGKBX
   allocationqHKCX   allowqIKDX   allyqJKEX   almostqKKFX   aloneqLKGX   alternativeqMKHX   amazingqNKIX
   ambassadorqOKJX	   ambulanceqPKKX   amendqQKLX   americasqRKMX   amputeeqSKNX   analystqTKOX   angerqUKPX   anglerqVKQX   angryqWKRX   animalqXKSX   announceqYKTX   announcementqZKUX   annualq[KVX   annuallyq\KWX   answerq]KXX   apartq^KYX	   apartmentq_KZX	   apologiseq`K[X   appealqaK\X   applaudqbK]X   applicationqcK^X   applyqdK_X   appointqeK`X   appointmentqfKaX   approachqgKbX   approvalqhKcX   approveqiKdX   aquaticqjKeX   archaeologicalqkKfX   areaqlKgX   argueqmKhX   ariseqnKiX   armedqoKjX   arrestqpKkX   arriveqqKlX   arrowqrKmX   arsenalqsKnX   arsonistqtKoX   arterialquKpX	   artilleryqvKqX   asbestosqwKrX   asideqxKsX   askqyKtX   assassinateqzKuX   assaultq{KvX   assessq|KwX
   assessmentq}KxX   assetq~KyX   assistqKzX
   assistanceq�K{X	   assuranceq�K|X
   astronomerq�K}X   asylumq�K~X   athleteq�KX   atrocityq�K�X   attackq�K�X   attemptq�K�X   attendq�K�X	   attendantq�K�X	   attentionq�K�X   attitudeq�K�X
   attractionq�K�X   auctionq�K�X   auditq�K�X   aussieq�K�X	   australiaq�K�X
   australianq�K�X	   authorityq�K�X	   availableq�K�X   avoidq�K�X   awaitq�K�X   awardq�K�X	   awarenessq�K�X   aynaouiq�K�X   backq�K�X   backingq�K�X   badlyq�K�X   baffleq�K�X   baftaq�K�X
   bairnsdaleq�K�X   baitq�K�X   balconyq�K�X   ballotq�K�X   banq�K�X
   bangladeshq�K�X   bankingq�K�X	   bankstownq�K�X   barrierq�K�X   baseq�K�X   bashq�K�X   basicq�K�X   basinq�K�X   basisq�K�X   battleq�K�X   bayernq�K�X   beachq�K�X   beatq�K�X   becomeq�K�X   bedouinq�K�X   beetleq�K�X   beginq�K�X   belgianq�K�X   believeq�K�X   believerq�K�X	   benchmarkq�K�X   benefitq�K�X   berthsq�K�X   betq�K�X   biddingq�K�X   bigq�K�X   billingq�K�X
   biologicalq�K�X   birthq�K�X   birthdayq�K�X   blackq�K�X   blameq�K�X   blastq�K�X   blatantq�K�X   blazeq�K�X   blazingq�K�X   blockq�K�X   bloodq�K�X   blueq�K�X   boardq�K�X   boardingq�K�X   bodyq�K�X   boggeq�K�X   bombq�K�X   bombardmentq�K�X   bombayq�K�X   bomberq�K�X   bombingq�K�X   bookieq�K�X   bookletq�K�X   boostq�K�X   borderq�K�X   bosnianq�K�X   bottleq�K�X   bottomq�K�X   bounceq�K�X   bowlerq�K�X   boxq�K�X	   boyfriendq�K�X   braveq�K�X   breakq�K�X   breakingq�K�X   breakoutq�K�X   breastq�K�X   breaststrokeq�K�X   bridgeq�K�X   bringq�K�X   britq�K�X   britishq�K�X	   broadcastq�K�X   broadcasterq�K�X   brokenq�K�X   brothelq�K�X   brotherq�K�X   brutalq�K�X   budgetq�K�X   buildq�K�X   builderq�K�X   buildingq�K�X   bullq�K�X   bulletq�K�X   bullyq�K�X   bullyingq�K�X
   bundesligaq�K�X   buoyantq�K�X   burdenq�K�X   burglaryq�K�X   burnq�K�X   burningq�K�X   buryq�K�X   bushfireq�K�X
   bushrangerq�K�X   businessq�K�X	   businesser   K�X   buyr  K�X   buyerr  K�X   bypassr  K�X   cabinetr  K�X   cadellr  M X   callr  MX	   caloundrar  MX	   cameramanr  MX   campaignr	  MX   canr
  MX   cancelr  MX   cancerr  MX	   candidater  MX   caner  M	X   cannabisr  M
X   cannonr  MX   canvassr  MX   canyonr  MX
   capabilityr  MX   capitalr  MX
   capitaliser  MX   captainr  MX   capturer  MX   caratr  MX   cardr  MX   cardiacr  MX   careerr  MX   carerr  MX
   caricaturer  MX   carryr  MX   caser  MX   casualtyr   MX   catchr!  MX   cattler"  MX   causer#  MX   cautionr$  MX   cautiousr%  M X   caver&  M!X	   celebrater'  M"X   celticr(  M#X
   censorshipr)  M$X   centr*  M%X   centralr+  M&X   centrer,  M'X   ceremonyr-  M(X   certainr.  M)X	   certaintyr/  M*X   cessnockr0  M+X   chairr1  M,X   chairmanr2  M-X	   challenger3  M.X   chamberr4  M/X   champr5  M0X   championr6  M1X   championshipr7  M2X   changer8  M3X   charader9  M4X   charger:  M5X   charterr;  M6X   chaser<  M7X
   checkpointr=  M8X   cheeser>  M9X   chelar?  M:X   chemicalr@  M;X   chickenrA  M<X   chiefrB  M=X   childrC  M>X	   childcarerD  M?X	   childhoodrE  M@X   childrenrF  MAX   chineserG  MBX   chokerH  MCX   chooserI  MDX   churchrJ  MEX   citizenrK  MFX   civilrL  MGX   civilianrM  MHX   claimrN  MIX   clashrO  MJX   classrP  MKX   cleanrQ  MLX   clearrR  MMX	   clearancerS  MNX   clearingrT  MOX   clemencyrU  MPX   clericrV  MQX   climbrW  MRX   clinicrX  MSX   cliprY  MTX   closerZ  MUX   closingr[  MVX   closurer\  MWX   cloudr]  MXX   clubr^  MYX   coachr_  MZX	   coalitionr`  M[X   coastra  M\X   coastalrb  M]X   cobawrc  M^X   cohesionrd  M_X   collaborationre  M`X   collapserf  MaX	   colleaguerg  MbX   colonialrh  McX   comeri  MdX   comebackrj  MeX	   commanderrk  MfX   commendrl  MgX   commentrm  MhX
   commissionrn  MiX   commitro  MjX
   commitmentrp  MkX   commonrq  MlX	   communityrr  MmX   companyrs  MnX
   compassionrt  MoX   competitionru  MpX	   complaintrv  MqX   completerw  MrX   complexrx  MsX   compoundry  MtX
   compromiserz  MuX   computerr{  MvX   concealr|  MwX   conceiver}  MxX   concernr~  MyX	   concernedr  MzX   concertr�  M{X   condemnr�  M|X	   conditionr�  M}X
   condolencer�  M~X   conductr�  MX
   confidencer�  M�X	   confidentr�  M�X   confirmr�  M�X   conflictr�  M�X   confrontr�  M�X	   confusionr�  M�X   congratulater�  M�X
   consciencer�  M�X   consentr�  M�X   consequencer�  M�X   conservationr�  M�X   conservativer�  M�X   considerr�  M�X   consolidater�  M�X   constructionr�  M�X   consultationr�  M�X   contactr�  M�X
   contagiousr�  M�X   containr�  M�X   containmentr�  M�X   contaminationr�  M�X   contestr�  M�X   contingencyr�  M�X   continuer�  M�X	   continuedr�  M�X   contractr�  M�X   contributionr�  M�X   controlr�  M�X   convictr�  M�X
   convictionr�  M�X   convoyr�  M�X   cooperationr�  M�X   coronerr�  M�X
   corruptionr�  M�X	   cosmonautr�  M�X   cossackr�  M�X   costr�  M�X   costlyr�  M�X   cottager�  M�X   cottonr�  M�X   couldr�  M�X   councilr�  M�X
   councillorr�  M�X   countr�  M�X   countryr�  M�X   coupler�  M�X   courser�  M�X   courtr�  M�X
   courthouser�  M�X   coverr�  M�X   coverager�  M�X   crackr�  M�X   craftr�  M�X	   craftsmenr�  M�X   crashr�  M�X   crazer�  M�X   creamr�  M�X   creanr�  M�X   creater�  M�X   creatorr�  M�X   credibilityr�  M�X   creditr�  M�X   crewr�  M�X   cricketr�  M�X	   cricketerr�  M�X   crimer�  M�X   criminalr�  M�X   crisisr�  M�X   criticr�  M�X   criticalr�  M�X	   criticiser�  M�X	   criticismr�  M�X   croonr�  M�X   cropr�  M�X   crossr�  M�X   crowr�  M�X   crownr�  M�X   cruder�  M�X   crueltyr�  M�X   cruiser�  M�X   crushr�  M�X   cryr�  M�X   cullr�  M�X   custodyr�  M�X   cutr�  M�X   cwealthr�  M�X   cycler�  M�X   damager�  M�X   dampenr�  M�X   dangler�  M�X   dater�  M�X   daubr�  M�X   daughterr�  M�X   deadliner�  M�X   deadlockr�  M�X   deadlyr�  M�X   dealr�  M�X   deathr�  M�X   debater�  M�X   decider�  M�X   decisionr�  M�X   declarer�  M�X   decliner�  M�X   dedicater�  M�X   deemr�  M�X   defeatr�  M�X   defectr�  M�X   defencer�  M�X   defendr�  M�X	   defensiver�  M�X   deficitr�  M�X   defraudr�  M�X   delayr�  M�X
   delegationr�  M�X   delightr�  M�X   deliverr�  M�X   demandr�  M�X   demolishr�  M�X	   demolisher�  M�X
   demolitionr�  M�X   demonr�  M�X   denguer�  M�X   dengue_outbreakr�  M�X   dentr   M�X   dentalr  M�X   denyr  M�X   departr  M�X	   departurer  M�X   deportr  M X   depositr  MX   deputyr  MX   deregulationr  MX   desaillyr	  MX   desalinationr
  MX   describer  MX   desertr  MX   deserver  MX   designerr  M	X   desirer  M
X	   desperater  MX
   despondentr  MX   destroyr  MX   destructionr  MX   detailr  MX   detainr  MX   detaineer  MX	   detentionr  MX   deterr  MX	   determiner  MX   developr  MX	   developerr  MX   developmentr  MX   devicer  MX   devilr  MX   deviser  MX   dialysisr   MX   dier!  MX
   differencer"  MX   digr#  MX   dinosaurr$  MX   dioufr%  M X	   diplomacyr&  M!X   diplomatr'  M"X	   directionr(  M#X   directorr)  M$X
   disappointr*  M%X   disarmr+  M&X   disasterr,  M'X
   disclosurer-  M(X
   discourager.  M)X	   discoveryr/  M*X   discriminationr0  M+X   discussr1  M,X   discusser2  M-X
   discussionr3  M.X   diseaser4  M/X
   disguisingr5  M0X   disgustr6  M1X   disillusionmentr7  M2X	   dismantler8  M3X   dismissr9  M4X	   dismissalr:  M5X   disputer;  M6X	   dissidentr<  M7X   distressr=  M8X   distributionr>  M9X   disturbr?  M:X	   diversionr@  M;X   dividerA  M<X   divisionrB  M=X   divorcerC  M>X   dockrD  M?X   dockerrE  M@X   doctorrF  MAX   dodgerG  MBX   dodgyrH  MCX   dollarrI  MDX   dolphinrJ  MEX   domesticrK  MFX   domestic_violencerL  MGX   dominaterM  MHX   donaterN  MIX   donationrO  MJX   doomrP  MKX   doorrQ  MLX   doperR  MMX   doralrS  MNX   dortmundrT  MOX   doublerU  MPX   doubtrV  MQX   downrW  MRX   downerrX  MSX   downfallrY  MTX   downpourrZ  MUX   doyler[  MVX   dozenr\  MWX   draftr]  MXX   drainr^  MYX   drainager_  MZX   draperr`  M[X   drawra  M\X   dreamrb  M]X   dredgerc  M^X   drenchrd  M_X   driftre  M`X   drillingrf  MaX   drinkrg  MbX   driverh  McX   driverri  MdX   dronerj  MeX   droprk  MfX   droughtrl  MgX   drownrm  MhX   drugrn  MiX   dryro  MjX   drylandrp  MkX   dukerq  MlX
   dumbledorerr  MmX   dumprs  MnX   dutchrt  MoX   eagerru  MpX   eaglerv  MqX   earlyrw  MrX   earnrx  MsX   earnerry  MtX   earthrz  MuX
   earthquaker{  MvX   easer|  MwX   easterr}  MxX   economicr~  MyX	   economistr  MzX   economyr�  M{X   edger�  M|X   editorr�  M}X	   educationr�  M~X   effectr�  MX   effluentr�  M�X   effortr�  M�X   egyptianr�  M�X   eighthr�  M�X   eldr�  M�X   elderlyr�  M�X   electr�  M�X   electionr�  M�X	   electoralr�  M�X   electricianr�  M�X   electricityr�  M�X
   electroluxr�  M�X   eligibler�  M�X	   eliminater�  M�X   emailr�  M�X   embassyr�  M�X   embedr�  M�X   embracer�  M�X   embryor�  M�X	   emergencyr�  M�X   emirater�  M�X   emissionr�  M�X	   emotionalr�  M�X   employeer�  M�X   employerr�  M�X
   employmentr�  M�X   enactr�  M�X	   encounterr�  M�X	   encourager�  M�X
   encouragedr�  M�X   endr�  M�X   endangerr�  M�X   endorsenentr�  M�X   enemyr�  M�X   engager�  M�X   enginer�  M�X   engineerr�  M�X   englandr�  M�X   englishr�  M�X   enoughr�  M�X   enqvistr�  M�X   enrager�  M�X   enrichr�  M�X   enriquer�  M�X   entallyr�  M�X   enterr�  M�X   entryr�  M�X   environmentr�  M�X   environmentalr�  M�X   envoyr�  M�X	   equaliserr�  M�X
   equestrianr�  M�X   eradicationr�  M�X   ergonr�  M�X   erosionr�  M�X   escaper�  M�X   escuder�  M�X   estater�  M�X   ethanolr�  M�X   ethicr�  M�X   ethnicr�  M�X   evacuater�  M�X   evaporationr�  M�X   eveningr�  M�X   eventr�  M�X   evidencer�  M�X   exactr�  M�X   examiner�  M�X   executer�  M�X	   executiver�  M�X   exhaustr�  M�X
   exhibitionr�  M�X   exiler�  M�X   expandr�  M�X	   expansionr�  M�X   expectr�  M�X   expectationr�  M�X	   expectingr�  M�X
   expeditionr�  M�X   expelr�  M�X   expenditurer�  M�X	   expensiver�  M�X
   experimentr�  M�X   experimentalr�  M�X   expertr�  M�X   explainr�  M�X   exploitationr�  M�X   explorationr�  M�X   explorer�  M�X	   explosionr�  M�X	   explosiver�  M�X   exportr�  M�X
   expressionr�  M�X	   expulsionr�  M�X   extendr�  M�X	   extensionr�  M�X   extrar�  M�X   extremer�  M�X	   extremismr�  M�X   eyer�  M�X   eyesorer�  M�X   facer�  M�X   facilityr�  M�X   factfiler�  M�X	   factionalr�  M�X   factor�  M�X   factorr�  M�X   factoryr�  M�X   fader�  M�X   failr�  M�X   fallr�  M�X   falloutr�  M�X   falser�  M�X   familyr�  M�X   farewellr�  M�X   farinasr�  M�X   farmr�  M�X   farmerr�  M�X   farmhandr�  M�X   fastr�  M�X   fatalr�  M�X   fatalityr�  M�X   fatherr�  M�X   favourr   M�X	   favouriter  M�X   fearr  M�X   featurer  M�X   federr  M�X   federalr  M X
   federationr  MX   federerr  MX   fedorovr  MX   feelr	  MX   femaler
  MX   fencer  MX   feralr  MX   fergier  MX   ferreror  M	X   ferryr  M
X   festivalr  MX   feverr  MX   fewr  MX	   feyenoordr  MX   fickler  MX   fieldr  MX   fiercer  MX   fifthr  MX   fightr  MX   fighterr  MX   fightingr  MX   figurer  MX   filer  MX   filmr  MX   finalr  MX   finalistr  MX   findr   MX   finer!  MX   finishr"  MX   finnishr#  MX   firer$  MX   fireballr%  M X   firefighterr&  M!X   firier'  M"X   firstr(  M#X   fisherr)  M$X	   fishermanr*  M%X   fisheryr+  M&X   fishingr,  M'X   flagr-  M(X   flamingor.  M)X   flashr/  M*X   fleer0  M+X   fleetr1  M,X   flemingr2  M-X   flightr3  M.X   flinderr4  M/X   floodr5  M0X   floodingr6  M1X   flowerr7  M2X   flyr8  M3X   focusr9  M4X   foldr:  M5X   followr;  M6X   footager<  M7X
   footballerr=  M8X   footingr>  M9X   footyr?  M:X   forbidr@  M;X   forcerA  M<X   forecastrB  M=X
   forecasterrC  M>X   foreignrD  M?X   forensicrE  M@X   foreseenrF  MAX   forestrG  MBX   forestryrH  MCX   forgetrI  MDX   forlanrJ  MEX   formrK  MFX   formalrL  MGX   formerrM  MHX   formularN  MIX   forumrO  MJX   forwardrP  MKX   fossilrQ  MLX   founderrR  MMX   fourthrS  MNX   foxrT  MOX   fragilerU  MPX   francerV  MQX   frankrW  MRX   fraudrX  MSX   freedomrY  MTX	   freestylerZ  MUX   freezer[  MVX   freezerr\  MWX   freightr]  MXX   frenchr^  MYX   freshr_  MZX   fridar`  M[X   friendlyra  M\X   frightenrb  M]X   frigorc  M^X   fruitrd  M_X   fruitpickerre  M`X
   frustratedrf  MaX   fundrg  MbX   fundingrh  McX   fundraisingri  MdX   funeralrj  MeX   futurerk  MfX   gainrl  MgX   galthierm  MhX   gambierrn  MiX   gamero  MjX   gangrp  MkX   gardenrq  MlX   gatecrasherrr  MmX   gatherrs  MnX   gearrt  MoX   gebrselassieru  MpX   gembrookrv  MqX   generalrw  MrX   geneticallyrx  MsX	   geraldtonry  MtX   germanrz  MuX   getr{  MvX   giantr|  MwX   giggsr}  MxX	   gilchristr~  MyX   giler  MzX	   gillespier�  M{X   gilmorer�  M|X   ginginr�  M}X	   gippslandr�  M~X   girdlerr�  MX   girlr�  M�X   giver�  M�X   glamourr�  M�X   globalr�  M�X   gloomr�  M�X   gloryr�  M�X   glover�  M�X   goallessr�  M�X   goldenr�  M�X	   goldfieldr�  M�X   golferr�  M�X   gonzalezr�  M�X
   governmentr�  M�X   governorr�  M�X   govtsr�  M�X   graderr�  M�X   grainr�  M�X   grandr�  M�X   grantr�  M�X   graper�  M�X   grazer�  M�X   grazierr�  M�X   greatr�  M�X   greecer�  M�X   greenr�  M�X   greener�  M�X
   greenpeacer�  M�X   grenader�  M�X   griffithr�  M�X   grosslyr�  M�X   groundr�  M�X   groundwaterr�  M�X   groupr�  M�X   growr�  M�X   growerr�  M�X   growthr�  M�X
   guantanamor�  M�X   guardr�  M�X   guerillar�  M�X	   guerrillar�  M�X   guider�  M�X   guiltyr�  M�X   gunr�  M�X   gunfirer�  M�X   gunmanr�  M�X   gunnedahr�  M�X   gunnerr�  M�X   gusmaor�  M�X   gutlessr�  M�X   gympier�  M�X
   gyrocopterr�  M�X   habitatr�  M�X   hackerr�  M�X
   hacktivistr�  M�X   hadjir�  M�X   hailr�  M�X	   hailstormr�  M�X	   hamackovar�  M�X   hancockr�  M�X   handr�  M�X   handler�  M�X   hangr�  M�X   happyr�  M�X   harmonyr�  M�X   harnessr�  M�X   harshr�  M�X   harvestr�  M�X   harveyr�  M�X   hatcheryr�  M�X   hater�  M�X   hawthornr�  M�X   haydenr�  M�X   headr�  M�X
   headmasterr�  M�X   healthr�  M�X   healthyr�  M�X   hearr�  M�X   hearingr�  M�X   heartr�  M�X
   heartbreakr�  M�X   heatr�  M�X   heatedr�  M�X   heavyr�  M�X   heavyweightr�  M�X   heftyr�  M�X   heightenr�  M�X
   helicopterr�  M�X   heninr�  M�X   henmanr�  M�X   henryr�  M�X   herbertr�  M�X   heritager�  M�X   heror�  M�X   herveyr�  M�X   hewittr�  M�X   hidder�  M�X   hider�  M�X   hidingr�  M�X	   highfieldr�  M�X
   highlanderr�  M�X	   highlightr�  M�X   highwayr�  M�X   hijackerr�  M�X   hikerr�  M�u(X	   hillgrover�  M�X	   hindrancer�  M�X   hintr�  M�X   hinzer�  M�X   historicr�  M�X
   historicalr�  M�X   historyr�  M�X   hitr�  M�X   hittingr�  M�X   hobartr�  M�X   hoddler�  M�X   hodger�  M�X   hodgsonr�  M�X   holdr�  M�X   holderr�  M�X   holer�  M�X   hollandr�  M�X   hollingworthr�  M�X   homer�  M�X   homelessr   M�X
   homosexualr  M�X   honourr  M�X   hooker  M�X   hooperr  M�X   hoper  M X   hopefulr  MX   horrorr  MX   horser  MX   hospicer	  MX   hospitalr
  MX   hospitaliser  MX   hospitalityr  MX   hostr  MX   hostager  M	X   hotelr  M
X   hotliner  MX   houllir  MX   houndr  MX   hourr  MX   houser  MX	   householdr  MX   housingr  MX   howardr  MX   huegillr  MX   humanr  MX   humanitarianr  MX   humanityr  MX   humphreyr  MX   hundredr  MX	   hungarianr  MX   hunterr  MX	   hurricaner   MX   hurtr!  MX   husbandr"  MX
   hystericalr#  MX   identifyr$  MX   identityr%  M X	   igelstromr&  M!X   illegalr'  M"X   illnessr(  M#X	   immediater)  M$X   immigrationr*  M%X
   immolationr+  M&X   immunisationr,  M'X   immuniser-  M(X   impactr.  M)X	   impactingr/  M*X
   impatiencer0  M+X   importr1  M,X   importationr2  M-X
   impoverishr3  M.X
   impressionr4  M/X   imprisonmentr5  M0X   improver6  M1X
   inadequater7  M2X
   inaugurater8  M3X	   incentiver9  M4X   incidentr:  M5X   includer;  M6X   incomer<  M7X   increaser=  M8X	   indemnityr>  M9X   independentr?  M:X   indexr@  M;X   indianrA  M<X
   indigenousrB  M=X
   indonesianrC  M>X   indoorrD  M?X   inductrE  M@X   indurainrF  MAX
   industrialrG  MBX   industryrH  MCX   infrastructurerI  MDX   injurerJ  MEX   injurierK  MFX   injuryrL  MGX   inmaterM  MHX   inquestrN  MIX   inquiryrO  MJX   insectrP  MKX   insistrQ  MLX
   inspectionrR  MMX	   inspectorrS  MNX   inspirerT  MOX   insteadrU  MPX   insultrV  MQX	   insurancerW  MRX   insurerrX  MSX   intenserY  MTX   interrZ  MUX   interestr[  MVX
   interestedr\  MWX   interimr]  MXX   internationalr^  MYX   internetr_  MZX	   interviewr`  M[X	   introducera  M\X   introductionrb  M]X   invaderc  M^X   invaderrd  M_X
   invalidatere  M`X   invasionrf  MaX   investigaterg  MbX   investigationrh  McX   investigatorri  MdX
   investmentrj  MeX   investorrk  MfX   inviterl  MgX   iranianrm  MhX   iraqirn  MiX   iraqisro  MjX   iraqsrp  MkX   irelandrq  MlX   irishrr  MmX
   irrigationrs  MnX	   irrigatorrt  MoX   irympleru  MpX   islamicrv  MqX   islamistrw  MrX   islandrx  MsX   islanderry  MtX   isolaterz  MuX   israelr{  MvX   israelir|  MwX   issuer}  MxX   italianr~  MyX   jailr  MzX	   jailhouser�  M{X   japanr�  M|X   japaneser�  M}X   jeremier�  M~X   jewellerr�  MX   jewishr�  M�X   jewistr�  M�X   jiranekr�  M�X   joblessr�  M�X   joeyr�  M�X   joinr�  M�X   jointr�  M�X   jooser�  M�X
   journalistr�  M�X   jubilantr�  M�X   judger�  M�X   judicialr�  M�X   jumpr�  M�X   jupiterr�  M�X   justicer�  M�X   juveniler�  M�X   kaiserslauternr�  M�X   kanimblar�  M�X   kayakerr�  M�X   keaner�  M�X   keater�  M�X   keelr�  M�X   keepr�  M�X   keppelr�  M�X   kesslerr�  M�X   kidnapr�  M�X   kidneyr�  M�X   killr�  M�X   kingr�  M�X   knifer�  M�X   knightr�  M�X   koreanr�  M�X
   kosciuszkor�  M�X   krogerr�  M�X   kuertenr�  M�X   kurdishr�  M�X   kuwaitr�  M�X   labelr�  M�X   laborr�  M�X   labourr�  M�X   ladyr�  M�X   laker�  M�X   lamentr�  M�X   landr�  M�X
   landholderr�  M�X   landingr�  M�X	   landslider�  M�X   langmackr�  M�X   larger�  M�X   lastr�  M�X   later�  M�X   laterr�  M�X   laughr�  M�X   launchr�  M�X   lavenderr�  M�X   lawyerr�  M�X   leadr�  M�X   leaderr�  M�X
   leadershipr�  M�X   leaguer�  M�X   learnr�  M�X   learnerr�  M�X   leaser�  M�X   leastr�  M�X   leaver�  M�X   lecturerr�  M�X   leedr�  M�X   legalr�  M�X   legislativer�  M�X	   leicesterr�  M�X   leiselr�  M�X   lengthr�  M�X   lentonr�  M�X   leopardr�  M�X   lesbianr�  M�X   lesterr�  M�X   lethalr�  M�X   letterr�  M�X   levelr�  M�X	   liabilityr�  M�X   liberalr�  M�X
   liberationr�  M�X   libertadorer�  M�X   libraryr�  M�X   licencer�  M�X   licenser�  M�X   lickr�  M�X	   lickliterr�  M�X   lier�  M�X   lifeliner�  M�X   lifesaver�  M�X	   lifesaverr�  M�X   lightr�  M�X	   lightningr�  M�X   lihirr�  M�X   likelyr�  M�X	   limestoner�  M�X   limitr�  M�X   liner�  M�X   linkr�  M�X   lionr�  M�X
   liquidatorr�  M�X   liquorr�  M�X   lismorer�  M�X   listr�  M�X   littler�  M�X	   liverpoolr�  M�X	   livestockr�  M�X   lobbyr�  M�X   lobsterr�  M�X   localr�  M�X   locallyr�  M�X   locustr�  M�X   logr�  M�X   loggerr�  M�X   lollyr�  M�X   longr�  M�X	   longreachr�  M�X   lookr�  M�X   loomr�  M�X   looser�  M�X   lootr�  M�X   loser�  M�X   lossr   M�X   lover  M�X
   lovenkrandr  M�X   lowr  M�X   lurr  M�X   lurkr  M X   madeirar  MX   majorr  MX   majorityr  MX   maker	  MX   makerr
  MX	   malaysianr  MX
   managementr  MX   managerr  MX   manufacturerr  M	X   manusr  M
X   marathonr  MX   marcher  MX   marginalr  MX   markr  MX   marketr  MX   marriager  MX	   martyrdomr  MX   massiver  MX   masterr  MX   matchr  MX	   maternityr  MX   matterr  MX   mayorr  MX   mayoralr  MX   mcdonaldr  MX   meanr  MX   measurer   MX
   meatworkerr!  MX   medalr"  MX   medicalr#  MX   mediciner$  MX   mediumr%  M X   meetr&  M!X   meetingr'  M"X	   melbourner(  M#X   memberr)  M$X
   membershipr*  M%X	   memorabler+  M&X   meningococcalr,  M'X   mentalr-  M(X   mentallyr.  M)X   merger/  M*X   mergerr0  M+X   messager1  M,X   metalr2  M-X   mexicanr3  M.X   meyerr4  M/X   militantr5  M0X   militaryr6  M1X   millr7  M2X   millionr8  M3X
   mindednessr9  M4X   minerr:  M5X   minimumr;  M6X   miningr<  M7X   ministerr=  M8X   ministryr>  M9X   minorr?  M:X   minuter@  M;X   mirerA  M<X   mishaprB  M=X   missrC  M>X   missilerD  M?X   missionrE  M@X   mobilerF  MAX   modifyrG  MBX   monarorH  MCX   moneyrI  MDX   monitorrJ  MEX   monthrK  MFX   monthlyrL  MGX   moralrM  MHX   morguerN  MIX   moroccanrO  MJX   mortgagerP  MKX   mosquerQ  MLX   motionrR  MMX
   motorcyclerS  MNX   motoristrT  MOX   mournrU  MPX   moverV  MQX   mudsliderW  MRX   mullrX  MSX   mummificationrY  MTX   murderrZ  MUX   murdererr[  MVX   musicr\  MWX   muzzler]  MXX   mysteryr^  MYX   nabr_  MZX   naiver`  M[X   namera  M\X   nasiriyarb  M]X	   nasiriyahrc  M^X   nationrd  M_X   nationalre  M`X   nativerf  MaX   naturalrg  MbX   naururh  McX   nearri  MdX   nearlyrj  MeX   needrk  MfX   neededrl  MgX   negativerm  MhX   neglectrn  MiX	   neighbourro  MjX   networkrp  MkX   newcomerrq  MlX	   newspaperrr  MmX   newspollrs  MnX   nigerianrt  MoX   nightru  MpX   ninthrv  MqX   noiserw  MrX   nominaterx  MsX   northry  MtX   northernrz  MuX   nuclearr{  MvX   numberr|  MwX   nurser}  MxX   nurseryr~  MyX   nursingr  MzX   obstructr�  M{X   occupyr�  M|X   offencer�  M}X   offenderr�  M~X   offerr�  MX   officerr�  M�X   officialr�  M�X   offsetr�  M�X   oldr�  M�X   olearyr�  M�X   oliver�  M�X   olympicr�  M�X   omaghr�  M�X   oncologyr�  M�X   openr�  M�X   openerr�  M�X	   operationr�  M�X   opponentr�  M�X   opposer�  M�X   opposedr�  M�X
   oppositionr�  M�X   optionr�  M�X   orderr�  M�X   oscarr�  M�X   oustr�  M�X   outdoorr�  M�X   outgoingr�  M�X   outlastr�  M�X   outlookr�  M�X   outskirtr�  M�X
   outstationr�  M�X   overr�  M�X	   overboardr�  M�X   overcomer�  M�X   overhaulr�  M�X   overheadr�  M�X   overtimer�  M�X   ownerr�  M�X   packager�  M�X   palacer�  M�X   palestinianr�  M�X   panelr�  M�X   panicr�  M�X   paperr�  M�X   parader�  M�X   parentr�  M�X
   parliamentr�  M�X   partialr�  M�X	   partiallyr�  M�X   partnerr�  M�X   partyr�  M�X   passr�  M�X	   passengerr�  M�X   pastoralr�  M�X   pathwayr�  M�X   patientr�  M�X   paymentr�  M�X   peacer�  M�X   peacefulr�  M�X   penaltyr�  M�X   penrithr�  M�X   peopler�  M�X   percentr�  M�X
   percentager�  M�X   perfectr�  M�X   perthr�  M�X   petrolr�  M�X   petrol_pricesr�  M�X   philippoussisr�  M�X   phoner�  M�X   pickr�  M�X
   pilgrimager�  M�X   pilotr�  M�X   pinr�  M�X   placer�  M�X   plaguer�  M�X   planr�  M�X   planer�  M�X   planningr�  M�X   plantr�  M�X   plantingr�  M�X   platformr�  M�X   playr�  M�X   playerr�  M�X   playingr�  M�X   pleadr�  M�X   pleaser�  M�X   pledger�  M�X   plummetr�  M�X	   pneumoniar�  M�X   pointr�  M�X   poisonr�  M�X	   poisoningr�  M�X   policer�  M�X	   policemanr�  M�X   policyr�  M�X   politicr�  M�X	   politicalr�  M�X
   politicianr�  M�X   pollr�  M�X   pollingr�  M�X   polluterr�  M�X	   pollutionr�  M�X   ponter�  M�X   ponyr�  M�X   poolr�  M�X   poorr�  M�X   poorlyr�  M�X
   populationr�  M�X   portr�  M�X   poser�  M�X   positionr�  M�X   positiver�  M�X   possibler�  M�X   postr�  M�X   postponer�  M�X	   potentialr�  M�X   potterr�  M�X   povertyr�  M�X   powerr�  M�X   poweredr�  M�X   praiser�  M�X   prayerr�  M�X   predictr�  M�X
   predictionr�  M�X
   preferencer�  M�X   pregnantr�  M�X   premierr�  M�X   premier_leaguer   M�X   premierer  M�X   premiershipr  M�X   premiumr  M�X   preparationr  M�X   preparer  M X   preparedr  MX   presencer  MX	   presidentr  MX   pressurer	  MX   pretextsr
  MX   previewr  MX   pricer  MX   primaryr  MX	   principler  M	X   priorityr  M
X   prisonr  MX   prisonerr  MX   privater  MX   privatisationr  MX	   privileger  MX   prober  MX   problemr  MX   processr  MX   producer  MX   producerr  MX
   productionr  MX   professionalr  MX   profiler  MX   profitr  MX   programr  MX   progressr  MX   projectr   MX   promiser!  MX   promoter"  MX   promptr#  MX
   propagandar$  MX   propertyr%  M X   proposalr&  M!X   prosecutionr'  M"X   prospectr(  M#X
   prosperityr)  M$X   protectr*  M%X
   protectionr+  M&X
   protectiver,  M'X   protestr-  M(X	   protesterr.  M)X   prover/  M*X   publicr0  M+X   publiclyr1  M,X   pullr2  M-X   punishr3  M.X
   punishmentr4  M/X   pushr5  M0X   qaedar6  M1X   quaker7  M2X	   qualifiedr8  M3X	   qualifierr9  M4X   qualifyr:  M5X   qualityr;  M6X
   quarantiner<  M7X   quarterr=  M8X   quashr>  M9X   queryr?  M:X   questionr@  M;X   quickrA  M<X	   quickfirerB  M=X   quitrC  M>X   quotarD  M?X   racerE  M@X   radiorF  MAX   radioactiverG  MBX   raidrH  MCX   rainrI  MDX   rainfallrJ  MEX   raiserK  MFX   rallyrL  MGX   rampagerM  MHX   ranchingrN  MIX   raperO  MJX   rarerP  MKX   raterQ  MLX	   ratepayerrR  MMX   reachrS  MNX   reactionrT  MOX   readrU  MPX   readyrV  MQX   realityrW  MRX
   reappointerX  MSX   reasonrY  MTX   rebuildrZ  MUX   recallr[  MVX   receiver\  MWX   recentr]  MXX   recklessr^  MYX	   recogniser_  MZX	   recommendr`  M[X   reconciliationra  M\X   recordrb  M]X   recoverrc  M^X   recoveryrd  M_X   recruitre  M`X	   recurrentrf  MaX   redbackrg  MbX   reducerh  McX	   reductionri  MdX
   redundancyrj  MeX   referrk  MfX   refereerl  MgX   reformrm  MhX	   reformistrn  MiX   refugeero  MjX   refusalrp  MkX   refuserq  MlX   regainrr  MmX   regattasrs  MnX   regimert  MoX   regionru  MpX   regionalrv  MqX   registerrw  MrX   regretrx  MsX   regularry  MtX	   regulatorrz  MuX   reintroducer{  MvX   rejectr|  MwX   relationshipr}  MxX   relaxr~  MyX   releaser  MzX   reliefr�  M{X   reliever�  M|X	   religiousr�  M}X   relocater�  M~X   relyr�  MX   remainr�  M�X
   remarkabler�  M�X   reminderr�  M�X   remover�  M�X   renalr�  M�X   reneger�  M�X   renewr�  M�X   reoffendr�  M�X   reopenr�  M�X   repairr�  M�X   repeatr�  M�X   replacer�  M�X   replacementr�  M�X   replayr�  M�X   reportr�  M�X
   reputationr�  M�X   requestr�  M�X   requirer�  M�X   rescuer�  M�X   researchr�  M�X
   researcherr�  M�X   reshaper�  M�X	   residencyr�  M�X   residentr�  M�X   residentialr�  M�X   resignr�  M�X   resistr�  M�X
   resistancer�  M�X
   resolutionr�  M�X   resolver�  M�X   resourcer�  M�X   responser�  M�X   responsibler�  M�X   restartr�  M�X   restockr�  M�X   restorationr�  M�X   restorer�  M�X   restrainr�  M�X	   restraintr�  M�X   restrictr�  M�X   restrictionr�  M�X   resultr�  M�X   resumer�  M�X   retailr�  M�X   retainr�  M�X   retaliationr�  M�X	   retentionr�  M�X   retirer�  M�X
   retirementr�  M�X   retracer�  M�X   retractr�  M�X   returnr�  M�X   reunionr�  M�X   reuniter�  M�X   revampr�  M�X   revealr�  M�X   revegetationr�  M�X   revenger�  M�X   reviewr�  M�X   reviser�  M�X   reviver�  M�X   revoltr�  M�X   rhoder�  M�X   rightr�  M�X   riser�  M�X   riskr�  M�X   rivalr�  M�X   roadr�  M�X   roadworkr�  M�X   robr�  M�X   robberr�  M�X   robbier�  M�X   rockr�  M�X   rocketr�  M�X   rompr�  M�X   rookier�  M�X   roper�  M�X   rotationr�  M�X   roundr�  M�X   router�  M�X   rowlingr�  M�X   ruler�  M�X   rulingr�  M�X   rumourr�  M�X   runr�  M�X   runningr�  M�X   ruralr�  M�X   russianr�  M�X   sackr�  M�X   safetyr�  M�X   saintr�  M�X   saler�  M�X   salinityr�  M�X   sanctionr�  M�X	   sandstormr�  M�X   sater�  M�X	   satelliter�  M�X	   satisfiedr�  M�X   satisfyr�  M�X   saver�  M�X   scallopr�  M�X   scarer�  M�X   scavenger�  M�X   scener�  M�X   scheduler�  M�X   schemer�  M�X   scholer�  M�X   schoolr�  M�X   schoolteacherr�  M�X   scorer�  M�X   scrapr�  M�X   scratchr�  M�X	   scrumbaser�  M�X   sculptorr�  M�X	   seachanger�  M�X   seafoodr�  M�X   sealr�  M�X   searchr�  M�X   seasonr�  M�X   seatr�  M�X   secondr�  M�X   secretr�  M�X   secretlyr�  M�X   sectionr   M�X   sectorr  M�X   securer  M�X   securityr  M�X   seedr  M�X   seekr  M X   seekerr  MX   seizer  MX	   selectionr  MX   sellr	  MX   sellerr
  MX   sendr  MX   sentencer  MX
   sentencingr  MX   separater  M	X   serbianr  M
X   seriesr  MX   seriousr  MX   server  MX   servicer  MX   setbackr  MX   settler  MX
   settlementr  MX   sevenr  MX   severalr  MX   sewerager  MX   shaker  MX   sharer  MX   shareholderr  MX   sharingr  MX   sharkr  MX   sharplyr  MX   shearr   MX   sheener!  MX   shelver"  MX   shieldr#  MX   shiner$  MX   shipr%  M X   shirer&  M!X   shirvor'  M"X   shockr(  M#X   shootr)  M$X   shoppingr*  M%X   shortr+  M&X   shortager,  M'X   showr-  M(X   showdownr.  M)X   shrugr/  M*X   shutr0  M+X	   sickeningr1  M,X   sider2  M-X   sideliner3  M.X   sieger4  M/X   sightr5  M0X   signr6  M1X   silencer7  M2X
   silverdomer8  M3X   simplyr9  M4X   singler:  M5X   sinkr;  M6X   sixr<  M7X   skater=  M8X   skateboardingr>  M9X   skillr?  M:X   skydiver@  M;X   slamrA  M<X   slashrB  M=X   slerC  M>X   slicerD  M?X   sliprE  M@X   slumprF  MAX   smallrG  MBX   smartrH  MCX   smelterrI  MDX   smokingrJ  MEX   smugglerK  MFX	   smugglingrL  MGX   snatchrM  MHX   sniffrN  MIX   soberrO  MJX   soccerrP  MKX   socialrQ  MLX   societyrR  MMX   solarrS  MNX   soldierrT  MOX   solemnrU  MPX   solutionrV  MQX   solverW  MRX   sourcerX  MSX   southrY  MTX   southernrZ  MUX   spacer[  MVX   sparkr\  MWX   speakr]  MXX   speakerr^  MYX   specialr_  MZX
   specialistr`  M[X   speciera  M\X   speedrb  M]X   speightrc  M^X   spillrd  M_X   splitre  M`X   spoilrf  MaX   sportrg  MbX   sportingrh  McX   spotri  MdX	   spotlightrj  MeX   sprayrk  MfX   spreadrl  MgX   sprinterrm  MhX   spurrn  MiX   spurtro  MjX   spyrp  MkX   squadrq  MlX   squarerr  MmX   squatterrs  MnX   stabrt  MoX   stabbingru  MpX   stackrv  MqX   staffrw  MrX   stafferrx  MsX   stagery  MtX   stallrz  MuX   stampr{  MvX   stancer|  MwX   starr}  MxX   startr~  MyX   starver  MzX   stater�  M{X	   statementr�  M|X   staticr�  M}X   stationr�  M~X	   statisticr�  MX   statusr�  M�X   stayr�  M�X   steadyr�  M�X   stealr�  M�X   steelr�  M�X   stickr�  M�X   stillr�  M�X   stockr�  M�X   stoddartr�  M�X   storager�  M�X   stormr�  M�X	   stragglerr�  M�X   straightr�  M�X   strandr�  M�X   strapr�  M�X	   strategicr�  M�X   strategyr�  M�X   strawr�  M�X   strayr�  M�X   streakr�  M�X
   strengthenr�  M�X   strickenr�  M�X   striker�  M�X   strikerr�  M�X   stroker�  M�X   strongr�  M�X   stronglyr�  M�X	   structurer�  M�X   struggler�  M�X   stuckr�  M�X   studentr�  M�X   studyr�  M�X   stumbler�  M�X   stunr�  M�X   stutterr�  M�X   subdivisionr�  M�X   subduer�  M�X
   submissionr�  M�X   subsidyr�  M�X   subwayr�  M�X   successr�  M�X
   successiver�  M�X   succumbsr�  M�X   suer�  M�X   sufferr�  M�X   sugarr�  M�X	   sugarcaner�  M�X   suicider�  M�X   suitr�  M�X   suitcaser�  M�X   summitr�  M�X   summonr�  M�X   superr�  M�X   superstitionr�  M�X   supplyr�  M�X   supportr�  M�X   surger�  M�X   surgeryr�  M�X   surplusr�  M�X   surpriser�  M�X	   surrenderr�  M�X   surveyr�  M�X   surviver�  M�X   survivorr�  M�X   suspectr�  M�X   suspendr�  M�X
   suspensionr�  M�X
   suspiciousr�  M�X   sustainabler�  M�X   swampr�  M�X   swanr�  M�X   swearr�  M�X   sweepr�  M�X	   sweetenerr�  M�X   swiftr�  M�X   swimmingr�  M�X   swindler�  M�X   swingr�  M�X   sydneyr�  M�X   symondr�  M�u(X   sympathyr�  M�X   syrianr�  M�X   syringer�  M�X   systemr�  M�X   tabler�  M�X   tacticr�  M�X   tagr�  M�X   taker�  M�X   takeoverr�  M�X   talkr�  M�X   tamer�  M�X   tankr�  M�X   targetr�  M�X	   tasmanianr�  M�X   taufelr�  M�X   teacherr�  M�X   teamr�  M�X   teenager�  M�X
   televisionr�  M�X   tellr�  M�X   tellerr�  M�X   temptr�  M�X   tenderr�  M�X   termr�  M�X	   territoryr�  M�X   terrorr�  M�X	   terrorismr�  M�X   testr�  M�X   testifyr�  M�X   textiler�  M�X   thailandr�  M�X   thankr�  M�X   theftr�  M�X   thiefr�  M�X   thinkr�  M�X   thirdr�  M�X   thorper�  M�X   thousandr�  M�X   thrashr�  M�X   threatr�  M�X   threatenr�  M�X   thrillerr�  M�X   throwr�  M�X   thumbr   M�X   thumpr  M�X   ticketr  M�X   tigerr  M�X   tightr  M�X
   tightlipper  M X   tikolor  MX   timberr  MX   timorr  MX   timoreser	  MX   tipr
  MX   tiredr  MX   tirrenor  MX   titler  MX   toastr  M	X   tobaccor  M
X   todayr  MX   toddlerr  MX   tomorrowr  MX   tonightr  MX   toolr  MX   toothr  MX   torrer  MX   torturer  MX   totalr  MX   touchr  MX   toughr  MX   tourr  MX   tourismr  MX   touristr  MX
   tournamentr  MX   towr  MX   townr   MX   townshipr!  MX   tracer"  MX   trackr#  MX   trader$  MX   tradingr%  M X	   traditionr&  M!X   traditionalr'  M"X
   traffickerr(  M#X   tragicr)  M$X   trailr*  M%X   trainr+  M&X   trainingr,  M'X	   transportr-  M(X   transsexualr.  M)X   travelr/  M*X   travir0  M+X   treasonr1  M,X   treasurer2  M-X	   treasurerr3  M.X	   treatmentr4  M/X   treatyr5  M0X   trebler6  M1X   trenchr7  M2X   trialr8  M3X   triangler9  M4X
   triathleter:  M5X   tributer;  M6X   trickr<  M7X   triggerr=  M8X   trimbler>  M9X   tripler?  M:X   triumphr@  M;X   trooprA  M<X   trophyrB  M=X   troubledrC  M>X   truancyrD  M?X   truckrE  M@X   trustrF  MAX   tryrG  MBX   tumutrH  MCX   tunnelrI  MDX
   turbulencerJ  MEX   turnrK  MFX   turnoutrL  MGX   tuskrM  MHX   tyrerN  MIX   umpiringrO  MJX   unbornrP  MKX	   uncertainrQ  MLX	   unchangedrR  MMX   unclearrS  MNX   unconcernedrT  MOX   undergoerU  MPX   underwayrV  MQX   unemploymentrW  MRX
   unexpectedrX  MSX   unfairrY  MTX   unfurlrZ  MUX   unhappyr[  MVX   unifyr\  MWX
   unilateralr]  MXX
   unimpresser^  MYX   unimpressedr_  MZX   uniter`  M[X   unitedra  M\X   unityrb  M]X   unknownrc  M^X   unlikelyrd  M_X   unmovere  M`X
   unoccupiedrf  MaX   unparalleledrg  MbX   unrestrh  McX   unswayeri  MdX   unveilrj  MeX   upbeatrk  MfX   upgraderl  MgX   upsetrm  MhX   uraniumrn  MiX   urgero  MjX   urgentrp  MkX   userrq  MlX   vaccinationrr  MmX   vacuumrs  MnX	   valuationrt  MoX   varietyru  MpX   vaultrv  MqX
   vegetationrw  MrX   venablerx  MsX   venuery  MtX   verdictrz  MuX   veteranr{  MvX	   viabilityr|  MwX   viabler}  MxX   victimr~  MyX	   victorianr  MzX   victoryr�  M{X   vigilantr�  M|X   villager�  M}X   violencer�  M~X   virusr�  MX   visitr�  M�X   voter�  M�X   voucherr�  M�X
   vulnerabler�  M�X   waitr�  M�X   waiver�  M�X   waler�  M�X
   walkinshawr�  M�X   walkoutr�  M�X   wanderr�  M�X   wantr�  M�X   warfarer�  M�X   warnr�  M�X   warningr�  M�X   washr�  M�X   wasimr�  M�X   waster�  M�X   watchr�  M�X   watchdogr�  M�X   watcherr�  M�X   waterr�  M�X   water_restrictionr�  M�X   water_supplyr�  M�X	   waterskier�  M�X   waughr�  M�X   waver�  M�X   wayner�  M�X   weaponr�  M�X   weatherr�  M�X   weekr�  M�X   weekendr�  M�X   welcomer�  M�X   welfarer�  M�X   wellr�  M�X   whaler�  M�X   wheatr�  M�X   whiner�  M�X   whiter�  M�X   whopperr�  M�X   wildcatr�  M�X
   wildernessr�  M�X   wilfulr�  M�X   willr�  M�X   winr�  M�X   windr�  M�X   windier�  M�X   winer�  M�X	   winegraper�  M�X	   winemakerr�  M�X   winlessr�  M�X   winnerr�  M�X   withdrawr�  M�X
   withdrawalr�  M�X	   withstandr�  M�X   witnessr�  M�X   wizardr�  M�X   wolfr�  M�X   womanr�  M�X   woodr�  M�X   woomerar�  M�X   workr�  M�X   workerr�  M�X   worldr�  M�X   wormr�  M�X   worryr�  M�X   worstr�  M�X   wouldr�  M�X   woundr�  M�X   woundedr�  M�X   wreakr�  M�X   writer�  M�X   wrongr�  M�X   yandinar�  M�X   yearr�  M�X	   yorkshirer�  M�X   youthr�  M�X   zoner�  M�X   abaloner�  M�X   abandonr�  M�X   abattoirr�  M�X   abider�  M�X
   aboriginalr�  M�X   abortionr�  M�X   abroadr�  M�X   absencer�  M�X   academicr�  M�X   acknowledger�  M�X   activer�  M�X   actorr�  M�X   administrationr�  M�X   adoptr�  M�X   advisoryr�  M�X   aerodynamicr�  M�X   agroundr�  M�X   aidr�  M�X   ailr�  M�X   algerianr�  M�X   americanr�  M�X   amoebar�  M�X   amputater�  M�X   anniversaryr�  M�X   anthraxr�  M�X   antidoter�  M�X   anwarr�  M�X   anxiousr�  M�X   appearr�  M�X   apprenticeshipr�  M�X   appropriater�  M�X   architecturalr�  M�X   armidaler�  M�X
   artificialr�  M�X   artificiallyr�  M�X   artistr�  M�X   aspirinr�  M�X   assassinationr�  M�X   assurer�  M�X   asthmar�  M�X   autopsyr�  M�X	   avalancher�  M�X   avertr�  M�X   babyr�  M�X	   babyholicr�  M�X   backlashr�  M�X
   backstroker 	  M�X   badr	  M�X   bananar	  M�X   basrar	  M�X   basslinkr	  M�X   battenr	  M 	X   beattier	  M	X   beggarr	  M	X   belittler	  M	X   bikier		  M	X   billionr
	  M	X   bindr	  M	X   biter	  M	X	   blackmailr	  M	X   blockader	  M		X	   bloodshedr	  M
	X   boatingr	  M	X   bolsterr	  M	X   bookr	  M	X   boomr	  M	X   borrowr	  M	X   bossr	  M	X   bowlingr	  M	X   bracer	  M	X   brainr	  M	X   braker	  M	X	   branchingr	  M	X   braveryr	  M	X   brawlr	  M	X   breachr	  M	X
   breastfeedr	  M	X   breedr	  M	X   briefr 	  M	X   brightr!	  M	X   brochurer"	  M	X   brumbier#	  M	X   bureaur$	  M	X
   bureaucratr%	  M 	X   burstr&	  M!	X
   bushwalkerr'	  M"	X   butcherr(	  M#	X	   butterflyr)	  M$	X   cainer*	  M%	X   calculationr+	  M&	X   callusr,	  M'	X   camerar-	  M(	X   campr.	  M)	X   campusr/	  M*	X   canadianr0	  M+	X   capacityr1	  M,	X   cappedr2	  M-	X   capsizer3	  M.	X
   careflightr4	  M/	X   carrierr5	  M0	X   castler6	  M1	X   casualr7	  M2	X	   catchmentr8	  M3	X   causingr9	  M4	X   ceaser:	  M5	X
   centraliser;	  M6	X	   centrebetr<	  M7	X
   challengerr=	  M8	X   chaosr>	  M9	X   chaplainr?	  M:	X   cheatr@	  M;	X   checkrA	  M<	X   cheerfulrB	  M=	X   chemistrC	  M>	X   chequerD	  M?	X   chillrE	  M@	X   chinarF	  MA	X   chiprG	  MB	X   choirrH	  MC	X   christchurchrI	  MD	X	   cigaretterJ	  ME	X   citerK	  MF	X   clarencerL	  MG	X   clarifyrM	  MH	X   cleaningrN	  MI	X   clijsterrO	  MJ	X   climaterP	  MK	X   clinchrQ	  ML	X   clonerR	  MM	X	   clubhouserS	  MN	X   clutchrT	  MO	X   coalminerU	  MP	X   coasterrV	  MQ	X   coffrW	  MR	X   colliderX	  MS	X	   collisionrY	  MT	X   colonrZ	  MU	X	   columnistr[	  MV	X   comedyr\	  MW	X   commemorater]	  MX	X   commerciallyr^	  MY	X   commissionerr_	  MZ	X   communicationr`	  M[	X   commuterra	  M\	X   companysrb	  M]	X
   comparablerc	  M^	X   competitivenessrd	  M_	X   complainre	  M`	X   comporf	  Ma	X   comraderg	  Mb	X   concederh	  Mc	X
   conferenceri	  Md	X   confusedrj	  Me	X
   connectionrk	  Mf	X   connollyrl	  Mg	X	   consulaterm	  Mh	X   consumerrn	  Mi	X	   contagionro	  Mj	X   contemptrp	  Mk	X
   contentionrq	  Ml	X
   contractorrr	  Mm	X
   contributers	  Mn	X   contributorrt	  Mo	X	   cooperateru	  Mp	X
   copenhagenrv	  Mq	X
   corinthianrw	  Mr	X	   corporaterx	  Ms	X   correspondentry	  Mt	X   cosgroverz	  Mu	X   costar{	  Mv	X
   counsellorr|	  Mw	X	   courtroomr}	  Mx	X   cowboyr~	  My	X	   crackdownr	  Mz	X   crankyr�	  M{	X   crayfishr�	  M|	X   creditorr�	  M}	X   creepr�	  M~	X
   criticallyr�	  M	X   crossbowr�	  M�	X   crosser�	  M�	X   crowdr�	  M�	X   crusaderr�	  M�	X   culturalr�	  M�	X   customr�	  M�	X   customerr�	  M�	X   cyanider�	  M�	X   cyberr�	  M�	X   cycloner�	  M�	X   cylinderr�	  M�	X   cypriotr�	  M�	X   dairyr�	  M�	X   darkenr�	  M�	X   darler�	  M�	X   davisr�	  M�	X   dealingr�	  M�	X   debitr�	  M�	X   debutr�	  M�	X   decapitationr�	  M�	X   deepenr�	  M�	X	   defaulterr�	  M�	X   defenderr�	  M�	X   defenser�	  M�	X   deferr�	  M�	X
   deliberater�	  M�	X   deliberatelyr�	  M�	X   denouncer�	  M�	X   densityr�	  M�	X   deployr�	  M�	X   deployedr�	  M�	X
   deploymentr�	  M�	X   derwentr�	  M�	X   destiner�	  M�	X	   devastater�	  M�	X	   dexterityr�	  M�	X   diabetesr�	  M�	X	   differentr�	  M�	X   diggerr�	  M�	X   dioxinr�	  M�	X
   diplomaticr�	  M�	X   directr�	  M�	X   disabledr�	  M�	X   disallowr�	  M�	X   disappearancer�	  M�	X
   discipliner�	  M�	X   discoverr�	  M�	X   dishr�	  M�	X   displayr�	  M�	X   disruptr�	  M�	X   dissolutionr�	  M�	X   disunityr�	  M�	X   diverser�	  M�	X	   diversityr�	  M�	X   dividedr�	  M�	X   djindjicr�	  M�	X   doggier�	  M�	X	   dominancer�	  M�	X	   downgrader�	  M�	X   dragonr�	  M�	X   dramaticr�	  M�	X   dredgingr�	  M�	X   easyr�	  M�	X	   economiser�	  M�	X   ectasyr�	  M�	X   edictr�	  M�	X   educatorr�	  M�	X   electrocuter�	  M�	X   eliminationr�	  M�	X   eliter�	  M�	X	   embarrassr�	  M�	X   emerger�	  M�	X   enforcer�	  M�	X
   engagementr�	  M�	X   enrolr�	  M�	X   ensurer�	  M�	X	   entertainr�	  M�	X   entirer�	  M�	X   entitlementr�	  M�	X
   entrapmentr�	  M�	X   environmentallyr�	  M�	X	   equipmentr�	  M�	X   eruptr�	  M�	X	   esperancer�	  M�	X   essayr�	  M�	X	   establishr�	  M�	X   esteemr�	  M�	X   eurobodallar�	  M�	X   europeanr�	  M�	X   excuser�	  M�	X	   executionr�	  M�	X   exemptr�	  M�	X	   exemptionr�	  M�	X   exerciser�	  M�	X   exodusr�	  M�	X   expenser�	  M�	X   exporterr�	  M�	X	   extraditer�	  M�	X	   extremistr�	  M�	X   extricationr�	  M�	X   facader�	  M�	X   factosr�	  M�	X   falterr�	  M�	X   fashionr�	  M�	X   fatiguer�	  M�	X   fatiguedr�	  M�	X   faultr�	  M�	X   feasibilityr�	  M�	X   featherr�	  M�	X   feelingr�	  M�	X   fiancer�	  M�	X   filthyr�	  M�	X   finaliser�	  M�	X   finallyr�	  M�	X   financer�	  M�	X	   financialr�	  M�	X   findingr�	  M�	X	   firebreakr�	  M�	X	   firefightr�	  M�	X
   firefighter�	  M�	X	   firepowerr�	  M�	X   fitnessr�	  M�	X   fixr�	  M�	X   flavellr 
  M�	X   flierr
  M�	X   flockr
  M�	X   flowr
  M�	X
   fluminenser
  M�	X   flutterr
  M 
X   footstepr
  M
X	   foreignerr
  M
X
   foreshadowr
  M
X   forger	
  M
X
   formidabler

  M
X   foyerr
  M
X   fracturer
  M
X   franticr
  M
X   freer
  M	
X   freelyr
  M

X   freewayr
  M
X	   fremantler
  M
X   friendr
  M
X   frogr
  M
X   frontr
  M
X	   furniturer
  M
X   gamblingr
  M
X
   gandolfinir
  M
X   generater
  M
X   ghanr
  M
X   gloomyr
  M
X   gor
  M
X   goalr
  M
X   governr
  M
X   gradr
  M
X	   grapeviner
  M
X
   greenhouser 
  M
X   greetr!
  M
X   gripr"
  M
X   grumbler#
  M
X   guestr$
  M
X	   guideliner%
  M 
X   hailedr&
  M!
X   haltr'
  M"
X   hamperr(
  M#
X   handsomer)
  M$
X   harbourr*
  M%
X   hardyr+
  M&
X	   harvesterr,
  M'
X
   harvestingr-
  M(
X   headhuntr.
  M)
X   heedr/
  M*
X   helenr0
  M+
X   helpr1
  M,
X   highr2
  M-
X	   hijackingr3
  M.
X   hirer4
  M/
X   holdingr5
  M0
X   holidayr6
  M1
X   homesicknessr7
  M2
X   hoodoor8
  M3
X   hostiler9
  M4
X   hotlyr:
  M5
X   hugher;
  M6
X   humbler<
  M7
X   hurdler=
  M8
X	   hypocrisyr>
  M9
X   ignorer?
  M:
X   imager@
  M;
X   imminentrA
  M<
X   imparjarB
  M=
X
   importancerC
  M>
X   imposerD
  M?
X
   impossiblerE
  M@
X   improvedrF
  MA
X   improvementrG
  MB
X	   inauguralrH
  MC
X   incenserI
  MD
X   inciterJ
  ME
X	   incursionrK
  MF
X   indecentrL
  MG
X   indiarM
  MH
X   indian_wellrN
  MI
X   indicaterO
  MJ
X   indierP
  MK
X   industrial_actionrQ
  ML
X
   inevitablerR
  MM
X   infantryrS
  MN
X	   infectionrT
  MO
X	   influencerU
  MP
X
   inhibitionrV
  MQ
X   injectrW
  MR
X   injuredrX
  MS
X   innerrY
  MT
X	   innisfailrZ
  MU
X   inputr[
  MV
X   instalr\
  MW
X   intelligencer]
  MX
X
   intensifier^
  MY
X   investr_
  MZ
X   invitationalr`
  M[
X   involvementra
  M\
X   iraqi_diplomatrb
  M]
X   ironmanrc
  M^
X	   irradiaterd
  M_
X   irreplaceablere
  M`
X   irreversiblerf
  Ma
X   itemrg
  Mb
X
   ivanisevicrh
  Mc
X   ivoryri
  Md
X   jacketrj
  Me
X   jayasuriyasrk
  Mf
X   jeerrl
  Mg
X   jitteryrm
  Mh
X   journeyrn
  Mi
X   justifyro
  Mj
X   kenyasrp
  Mk
X   kickrq
  Ml
X   killerrr
  Mm
X   killingrs
  Mn
X   kindredrt
  Mo
X   kittyru
  Mp
X	   klitschkorv
  Mq
X   knowrw
  Mr
X   lashrx
  Ms
X   leakry
  Mt
X   legalityrz
  Mu
X   lemonr{
  Mv
X   letr|
  Mw
X   liabler}
  Mx
X   licenseer~
  My
X   lifer
  Mz
X
   lifesavingr�
  M{
X   liftr�
  M|
X   lightingr�
  M}
X
   limitationr�
  M~
X   linerr�
  M
X   liquidr�
  M�
X   literacyr�
  M�
X   litrer�
  M�
X   liver�
  M�
X   lodger�
  M�
X   lookoutr�
  M�
X   lottor�
  M�
X   lowerr�
  M�
X   loyalistr�
  M�
X   loyaltyr�
  M�
X   lyrebirdr�
  M�
X   machiner�
  M�
X
   madagascarr�
  M�
X   magpier�
  M�
X   mailr�
  M�
X   maintainr�
  M�
X   manr�
  M�
X   mandater�
  M�
X   manlyr�
  M�
X   manslaughterr�
  M�
X   manualr�
  M�
X   marchr�
  M�
X   marillir�
  M�
X   mariner�
  M�
X   martinr�
  M�
X   martyrr�
  M�
X   maskr�
  M�
X   masser�
  M�
X
   mastermindr�
  M�
X   mater�
  M�
X   materialr�
  M�
X   mbekir�
  M�
X   mccainr�
  M�
X   mcewenr�
  M�
X   meltingr�
  M�
X   memorialr�
  M�
X   menacer�
  M�
X   menindeer�
  M�
X
   meningitisr�
  M�
X   methaner�
  M�
X   metrer�
  M�
X   micromanager�
  M�
X   middler�
  M�
X	   milosevicr�
  M�
X   minimalr�
  M�
X   minimiser�
  M�
X   miracler�
  M�
X
   misconductr�
  M�
X   misleadr�
  M�
X   misrepresentedr�
  M�
X   missingr�
  M�
X   missing_yachtsmanr�
  M�
X   mixr�
  M�
X   mixedr�
  M�
X   modelr�
  M�
X   momentumr�
  M�
X   monumentr�
  M�
X   moraler�
  M�
X
   moratoriumr�
  M�
X   mortarr�
  M�
X   motherr�
  M�
X   motivater�
  M�
X	   motorbiker�
  M�
X   mountr�
  M�
X   movementr�
  M�
X   mozzier�
  M�
X   mugaber�
  M�
X   musicalr�
  M�
X   muter�
  M�
X   narrowr�
  M�
X   neanderthalr�
  M�
X	   necessityr�
  M�
X   negotiationr�
  M�
X   neverr�
  M�
X   nordicr�
  M�
X   notchr�
  M�
X   obesityr�
  M�
X   observerr�
  M�
X   officer�
  M�
X   offshorer�
  M�
X   okayr�
  M�
X
   oncologistr�
  M�
X   ongoingr�
  M�
X   opalr�
  M�
X   operatorr�
  M�
X   orchidr�
  M�
X   orderlyr�
  M�
X	   organiserr�
  M�
X   outbreakr�
  M�
X   outburstr�
  M�
X   outdatedr�
  M�
X   outerr�
  M�
X   outlawr�
  M�
X   outliver�
  M�
X   outsider�
  M�
X   outsourcingr�
  M�
X   overallr�
  M�
X   overconfidencer�
  M�
X
   overflightr�
  M�
X	   overnightr�
  M�
X   overseasr�
  M�
X   overseer�
  M�
X   overturnr�
  M�
X   oxfamr�
  M�
X   oxygenr�
  M�
X   packr�
  M�
X   packerr�
  M�
X   packingr�
  M�
X
   paedophiler�
  M�
X   paintr�
  M�
X	   pakistanir�
  M�
X   pandar�
  M�
X	   parachuter�
  M�
X   parachutingr�
  M�
X   parentalr�
  M�
X   parliamentaryr�
  M�
X   partnershipr�
  M�
X   pasmincor�
  M�
X   passionr�
  M�
X   pastoralistr�
  M�
X   patchr�
  M�
X   patheticr�
  M�
X
   peacefullyr�
  M�
X   peacekeepingr   M�
X   peakr  M�
X   pelletr  M�
X   pennyr  M�
X   performr  M�
X	   permanentr  M X   personr  MX   personalr  MX   petitionr  MX   phantomr	  MX   phaser
  MX   photographyr  MX   piggeryr  MX   pilbarar  MX   pinchr  M	X   pipeliner  M
X   pitchr  MX   placingr  MX   plannerr  MX
   plantationr  MX   plasticr  MX   pleasedr  MX   plotr  MX   plunger  MX   poachr  MX   podiumr  MX   poetr  MX	   pointlessr  MX   poiser  MX   pokyr  MX   pollockr  MX   pompeyr  MX   ponderr   MX   pontingr!  MX   poppyr"  MX   popularr#  MX
   popularityr$  MX   possessr%  M X   possibilityr&  M!X   posthumouslyr'  M"X   poundr(  M#X   powderr)  M$X	   powerliner*  M%X   practicer+  M&X   practiser,  M'X   prayr-  M(X	   pregnancyr.  M)X   presentr/  M*X   presidentialr0  M+X	   pressuredr1  M,X   pretzelr2  M-X   prevailr3  M.X   preventr4  M/X
   preventionr5  M0X   previousr6  M1X   prizer7  M2X   progressingr8  M3X   prohibitr9  M4X   proposer:  M5X
   prosecutorr;  M6X   prostitutionr<  M7X   provider=  M8X   provocationr>  M9X   psychiatristr?  M:X   psychologistr@  M;X	   publicistrA  M<X   punchrB  M=X   pursuerC  M>X   pylonrD  M?X
   qualifyingrE  M@X   quieterrF  MAX   quollrG  MBX   rabbitrH  MCX   racialrI  MDX   racismrJ  MEX   racistrK  MFX   radicalrL  MGX   ragerM  MHX   raiderrN  MIX   rankrO  MJX   rankingrP  MKX   rapidrQ  MLX   rapistrR  MMX   ratfierS  MNX   rationrT  MOX   rattlerU  MPX   ravagerV  MQX   rebelrW  MRX	   recapturerX  MSX   recederY  MTX	   recessionrZ  MUX
   reconsiderr[  MVX   recorderr\  MWX
   recreationr]  MXX   redeployr^  MYX   redevelopmentr_  MZX   regardr`  M[X
   registeredra  M\X   rehabilitationrb  M]X   reinforcementrc  M^X   reinventrd  M_X   relatedre  M`X   relationrf  MaX   relativerg  MbX   relayrh  McX   relishri  MdX   rememberrj  MeX   renamerk  MfX   resignationrl  MgX   respectrm  MhX   respiratoryrn  MiX   responsibilityro  MjX
   responsiverp  MkX   restrq  MlX   restaterr  MmX
   restaurantrs  MnX   restaurateurrt  MoX   retailerru  MpX   rethinkrv  MqX   retreatrw  MrX   retrieverx  MsX
   revelationry  MtX   revenuerz  MuX   ribbonr{  MvX   rider|  MwX   riverr}  MxX	   riverlandr~  MyX   roarr  MzX   rollr�  M{X   ronaldor�  M|X   roofsr�  M}X   rooneyr�  M~X   roosterr�  MX   roughr�  M�X   roverr�  M�X   rowr�  M�X   rowingr�  M�X   royalr�  M�X   rudderr�  M�X   ruddockr�  M�X   rugbyr�  M�X   rumbler�  M�X   runawayr�  M�X   ryler�  M�X   saddamr�  M�X   safer�  M�X   sailingr�  M�X   sailorr�  M�X   saleyardr�  M�X   samoar�  M�X   samprasr�  M�X	   sanctuaryr�  M�X   sandr�  M�X
   sandalwoodr�  M�X   sanderr�  M�X
   sangakkarar�  M�X   saudir�  M�X   savager�  M�X   sawmillr�  M�X   scaler�  M�X   scandalr�  M�X   scather�  M�X   schnyderr�  M�X   schoolier�  M�X	   schoolingr�  M�X	   schroederr�  M�X   schwabr�  M�X   sciencer�  M�X	   scientistr�  M�X   scotr�  M�X   screenr�  M�X	   screeningr�  M�X   scrutinyr�  M�X   scullyr�  M�X	   sculpturer�  M�X   seagullr�  M�X   searcherr�  M�X   seekingr�  M�X   seizurer�  M�X   seler�  M�X   selectorr�  M�X   senatorr�  M�X   seniorr�  M�X	   sentimentr�  M�X
   separatistr�  M�X   sequinr�  M�X	   seriouslyr�  M�X   sessionr�  M�X   settingr�  M�u(X   seventhr�  M�X   severer�  M�X   sewager�  M�X   sexuallyr�  M�X   shackr�  M�X   shadowr�  M�X   share_marketr�  M�X   sharpenr�  M�X   shaughnessyr�  M�X   sheedyr�  M�X   sheepr�  M�X
   sheppartonr�  M�X
   shevchenkor�  M�X   shimanger�  M�X   shooterr�  M�X   shootingr�  M�X   shopr�  M�X   shopperr�  M�X   shortlyr�  M�X   shotr�  M�X   shouldr�  M�X   shoulderr�  M�X
   showgroundr�  M�X   showingr�  M�X   shunr�  M�X   shuttler�  M�X   siblingr�  M�X   signager�  M�X   signalr�  M�X   siliconr�  M�X   silverr�  M�X   simonir�  M�X   sisterr�  M�X   siter�  M�X   sizzlingr�  M�X   skaifer�  M�X   skaser�  M�X   skiingr�  M�X   skilledr�  M�X   skyr�  M�X   skywr�  M�X   slackr�  M�X   slainr�  M�X   slappingr�  M�X   slaterr�  M�X   slaver�  M�X   sleepr�  M�X   slider�  M�X   slipperyr�  M�X   slowr�  M�X   slowlyr�  M�X   smallerr�  M�X   smashr�  M�X   smellr�  M�X   smoker�  M�X   smugglerr�  M�X   snaker�  M�X   sniperr�  M�X   snowboarderr�  M�X   snowier�  M�X   snowtownr�  M�X	   socceroosr�  M�X
   softballerr�  M�X   solomonr�  M�X   solventr�  M�X   soorleyr�  M�X   sopranor�  M�X	   sorenstamr   M�X   sounessr  M�X   spanishr  M�X   specialisedr  M�X	   spectatorr  M�X   speculationr  M X   speechr  MX   spellr  MX   spendr  MX   spendingr	  MX   spiltr
  MX   spiritr  MX	   spokesmanr  MX   spreer  MX   sprinbokr  M	X
   springborgr  M
X	   sprinklerr  MX   spurnr  MX   spyingr  MX   squeezer  MX   stackerr  MX   staffingr  MX	   stalemater  MX   stalkr  MX   standr  MX   standardr  MX   starterr  MX   ster  MX   steerr  MX   stellarr  MX   stepr  MX   sterreyr  MX   stingerr   MX   stomachr!  MX   stompingr"  MX   stoner#  MX   stopr$  MX   stopoverr%  M X   strainr&  M!X   strawsr'  M"X   streetr(  M#X   strengthr)  M$X   strictr*  M%X   stripr+  M&X   stunningr,  M'X	   stuttgartr-  M(X   styler.  M)X   subjectr/  M*X
   substituter0  M+X
   subversiver1  M,X   suggestr2  M-X
   suggestionr3  M.X   sunracer4  M/X   sunriser5  M0X   supr6  M1X   supercomputerr7  M2X   supermarketr8  M3X   supplementaryr9  M4X	   supremacyr:  M5X   surfr;  M6X   surroundr<  M7X	   surveyingr=  M8X   survivalr>  M9X   svenr?  M:X   swainr@  M;X   swazirA  M<X   swimmerrB  M=X   swiperC  M>X   swissrD  M?X	   symposiumrE  M@X   symptomrF  MAX   szaborG  MBX	   tablelandrH  MCX   tabletrI  MDX   tacklerJ  MEX   tadpolerK  MFX   taipanrL  MGX   talentrM  MHX   tallisrN  MIX   tamworthrO  MJX   tanevularP  MKX   tangararQ  MLX   taperR  MMX   taperrS  MNX   tariffrT  MOX   tassierU  MPX   tavernrV  MQX	   technicalrW  MRX
   technologyrX  MSX   teenrY  MTX   teenagerrZ  MUX   telstrar[  MVX   tennantr\  MWX   tennisr]  MXX   tenser^  MYX   tensionr_  MZX   terminalr`  M[X	   terrifiedra  M\X	   terroristrb  M]X   testingrc  M^X   thankyourd  M_X   thighre  M`X	   threesomerf  MaX   thrillrg  MbX   thrustrh  McX   thunderbirdri  MdX   thunderstormrj  MeX   thwaiterk  MfX   tightenrl  MgX   timerm  MhX   timelyrn  MiX   tippedro  MjX   tissuerp  MkX   togetherrq  MlX	   tolerancerr  MmX   tongars  MnX	   toowoombart  MoX   topplingru  MpX   tortoiserv  MqX   tossrw  MrX   touchingrx  MsX   toxicry  MtX   toyworldrz  MuX   trafficr{  MvX   trailerr|  MwX   trainerr}  MxX   tranquiliserr~  MyX   transferr  MzX   transitr�  M{X   transparencyr�  M|X
   transplantr�  M}X	   traumaticr�  M~X
   traumatiser�  MX	   travellerr�  M�X   trawlerr�  M�X   treatr�  M�X   trefoilr�  M�X   tremorr�  M�X	   trezeguetr�  M�X   tribunalr�  M�X   trimr�  M�X   tropfr�  M�X   tropicalr�  M�X   troubler�  M�X   truckerr�  M�X   truckier�  M�X   truckingr�  M�X   tuckeyr�  M�X   tugboatr�  M�X   tumbler�  M�X   tupour�  M�X   turkeyr�  M�X   turkishr�  M�X   turnbullr�  M�X   turtler�  M�X   tweedr�  M�X   twelfthr�  M�X   tysonr�  M�X   ulirachr�  M�X   ulsterr�  M�X	   ultimatumr�  M�X
   ultralightr�  M�X   unbeatenr�  M�X   uncertaintyr�  M�X   undecider�  M�X	   undecidedr�  M�X   underager�  M�X
   undercoverr�  M�X   undergroundr�  M�X
   undeterredr�  M�X	   unethicalr�  M�X   unfitr�  M�X   unforgivabler�  M�X   unharmer�  M�X   unhookedr�  M�X   unicefr�  M�X   unionr�  M�X   unitr�  M�X
   unlicencedr�  M�X	   unsecuredr�  M�X   unsurer�  M�X   unusualr�  M�X   updater�  M�X   upgradedr�  M�X   upperr�  M�X   utahr�  M�X   vacciner�  M�X   vailer�  M�X   vandalr�  M�X	   vandalismr�  M�X   vanstoner�  M�X   vehicler�  M�X   venterr�  M�X   venturer�  M�X   venusr�  M�X   verificationr�  M�X
   verstappenr�  M�X   vialr�  M�X   victoriar�  M�X   videor�  M�X   vidukar�  M�X   vidukasr�  M�X   vieirar�  M�X   villagerr�  M�X   vintager�  M�X   violentr�  M�X   virginr�  M�X   virtualr�  M�X   visionr�  M�X   visitorr�  M�X   vitalr�  M�X	   voluntaryr�  M�X	   volunteerr�  M�X   voterr�  M�X   votingr�  M�X   vowler�  M�X   wager�  M�X   wagonr�  M�X   waitingr�  M�X   walesr�  M�X   walkr�  M�X   walkerr�  M�X   wallr�  M�X   wallabyr�  M�X   wallir�  M�X	   wanderingr�  M�X   waratahsr�  M�X   warhorser�  M�X   warner�  M�X   warplaner�  M�X   warriorr�  M�X   washingr�  M�X	   waterfallr�  M�X   waterwayr�  M�X   watkinr�  M�X   wedr�  M�X   weddingr�  M�X   weighr�  M�X   weightr�  M�X   wellmanr�  M�X	   wesfarmerr�  M�X   westernr�  M�X	   westernerr�  M�X   wetlandr�  M�X   whatmorer�  M�X   wheelr�  M�X   wicketr�  M�X   wicklowr�  M�X   widenr�  M�X   widner�  M�X   widowr�  M�X   wildlifer�  M�X
   williamsonr�  M�X   willingnessr�  M�X   wimmerar�  M�X   winchr�  M�X   wiper   M�X   wishr  M�X   womenr  M�X   woodchipr  M�X
   woolgrowerr  M�X	   woolworthr  M X   wordr  MX   workingr  MX   worksafer  MX	   worldwider	  MX   worser
  MX   wrangler  MX   wrapr  MX   wreckr  MX	   writedownr  M	X   writerr  M
X   yachtr  MX	   yachtsmanr  MX   yarakar  MX   yemenir  MX   youngr  MX	   youngsterr  MX   zabaletar  MX   abarer  MX   abdicater  MX   abductr  MX   ablazer  MX	   aboriginer  MX   abortr  MX	   abundancer  MX   accentr  MX   accountabilityr  MX
   accusationr   MX   achiever!  MX   achievementr"  MX   acquisitionr#  MX   acquitr$  MX   actr%  M X   addictr&  M!X	   addictionr'  M"X   adjustr(  M#X   adoptionr)  M$X   adultr*  M%X   advertisingr+  M&X
   aftershockr,  M'X   ager-  M(X   agfr.  M)X	   alcoholicr/  M*X   algaer0  M+X   alinghir1  M,X	   allegedlyr2  M-X   alsacer3  M.X   altercationr4  M/X	   aluminiumr5  M0X   ambitionr6  M1X	   ambitiousr7  M2X	   amendmentr8  M3X   ameryr9  M4X   aminor:  M5X
   ammunitionr;  M6X   amnestyr<  M7X   amrozir=  M8X	   ancestralr>  M9X   anchorr?  M:X   ancientr@  M;X   andersonrA  M<X   anglerB  M=X
   annihilaterC  M>X	   antarcticrD  M?X   anticrE  M@X   apparentrF  MAX   arabicrG  MBX   arafatrH  MCX   arbitrationrI  MDX
   arbitratorrJ  MEX   archaeologistrK  MFX	   architectrL  MGX	   argentinerM  MHX   argentinianrN  MIX   argumentrO  MJX   armourrP  MKX   arnhemrQ  MLX   arrangerR  MMX   arsonrS  MNX   arthurrT  MOX   artworkrU  MPX   asherV  MQX   asianrW  MRX   assassinrX  MSX	   assistantrY  MTX   athensrZ  MUX   athleticr[  MVX   atleticor\  MWX   atsicr]  MXX   austr^  MYX   austeelr_  MZX   autumnr`  M[X   aviationra  M\X	   avoidancerb  M]X   awarerc  M^X   bacherrd  M_X
   backpackerre  M`X	   backpedalrf  MaX   baghdadrg  MbX   balancerh  McX   ballackri  MdX   ballaratrj  MeX
   ballooningrk  MfX   bangladeshsrl  MgX   bankrm  MhX   baptistrn  MiX   bargainro  MjX
   bargainingrp  MkX   barginrq  MlX   barrichellorr  MmX   bartholomeuzrs  MnX   baseballrt  MoX	   batchelorru  MpX   batemanrv  MqX	   bathhouserw  MrX   baxterrx  MsX   bearry  MtX   beazleyrz  MuX	   beekeeperr{  MvX   behaver|  MwX   behindr}  MxX   belgiumr~  MyX   beller  MzX   belohvosciksr�  M{X   benchr�  M|X   bendigor�  M}X   bergerr�  M~X   bergkampr�  MX   bevanr�  M�X   bewarer�  M�X   biasedr�  M�X   bickerr�  M�X	   bickeringr�  M�X	   bilateralr�  M�X   bilbyr�  M�X   billionairer�  M�X	   biologistr�  M�X   birdr�  M�X   blackallr�  M�X   blackoutr�  M�X
   blackshirtr�  M�X   blaker�  M�X   bleedr�  M�X   blendr�  M�X   blighr�  M�X   blightr�  M�X   blindr�  M�X   blitzr�  M�X   bloker�  M�X   bloodierr�  M�X   bloodyr�  M�X
   boardshortr�  M�X   boatr�  M�X   boksicr�  M�X   bombardr�  M�X   bonlacr�  M�X   bonusr�  M�X   boomer�  M�X   botchr�  M�X   boulamir�  M�X   bourker�  M�X   brackr�  M�X   brackenr�  M�X   brandr�  M�X	   breakdownr�  M�X   breakthroughr�  M�X   breedingr�  M�X	   briefcaser�  M�X   brightenr�  M�X   brinkr�  M�X   britainr�  M�X   broadr�  M�X	   broadbandr�  M�X   brogdenr�  M�X   brokingr�  M�X   broncor�  M�X	   brookdaler�  M�X   broomer�  M�X   brownr�  M�X   brownlowr�  M�X   brundler�  M�X   bryantr�  M�X   bucherr�  M�X   buddhistr�  M�X   bulldogr�  M�X   bumperr�  M�X   bunnyr�  M�X   burier�  M�X   burker�  M�X   burmar�  M�X
   burrendongr�  M�X   busr�  M�X
   bushmasterr�  M�X   busterr�  M�X   butlerr�  M�X   buttonr�  M�X   caleyr�  M�X   callerir�  M�X   callousr�  M�X   cambodiar�  M�X	   cambodianr�  M�X   campaigningr�  M�X   camplinr�  M�X   cancellationr�  M�X   candleholderr�  M�X
   canegrowerr�  M�X   canoeistr�  M�X   canyonerr�  M�X   capabler�  M�X   capriatir�  M�X	   captaincyr�  M�X   captiver�  M�X   cardiologistr�  M�X   carewr�  M�X   carnager�  M�X   carparkr�  M�X   carpentariar�  M�X   carrr�  M�X
   carseldiner�  M�X   casinor�  M�X   cataractr�  M�X   categoryr�  M�X   catholicr�  M�X	   cattlemanr�  M�X   caucusr�  M�X   causedr�  M�X	   ceasefirer�  M�X   celebrationr�  M�X   celtr�  M�X   cemeteryr�  M�X   censorr�  M�X   censusr�  M�X
   centrelinkr�  M�X   centuryr�  M�X   cfmeur�  M�X   chainr�  M�X   chancer�  M�X   chaoticr�  M�X   chappellr�  M�X   charityr�  M�X   charlestownr�  M�X   cheapr�  M�X   cherryr�  M�X   chestr�  M�X   chewr�  M�X   chievor�  M�X   childcare_centrer�  M�X   chileanr�  M�X   choicer�  M�X   chromer�  M�X   chunkyr�  M�X   cityr   M�X   citylinkr  M�X   civicr  M�X   clamberr  M�X   clampr  M�X   clarkr  M X   clarker  MX   classicr  MX   classyr  MX   clotr	  MX
   clydesdaler
  MX	   coastliner  MX   coler  MX   collarr  MX   colleger  M	X   collinr  M
X	   collusionr  MX   colombiar  MX	   colombianr  MX	   columbianr  MX   combatr  MX   combiner  MX   comfortr  MX
   commercialr  MX   commericialr  MX	   committedr  MX   commonplacer  MX
   competencer  MX
   compliancer  MX
   compulsoryr  MX   concerns_airer  MX   concerns_airedr  MX   concorder   MX   condemnationr!  MX	   conductorr"  MX   confessr#  MX   confiner$  MX   confiscatedr%  M X   conscientiousr&  M!X   consistencyr'  M"X   consultr(  M#X
   consultantr)  M$X   contaminater*  M%X
   contingentr+  M&X   contriter,  M'X   controversialr-  M(X   converger.  M)X   coomar/  M*X	   copyrightr0  M+X   coralr1  M,X   corambar2  M-X   corinithianr3  M.X   corkr4  M/X
   coronationr5  M0X   coronialr6  M1X   corporationr7  M2X   correctionalr8  M3X   corserr9  M4X   cosmeticr:  M5X   cosmicr;  M6X   costellor<  M7X	   coulthardr=  M8X   counselr>  M9X   counsellingr?  M:X   counterattackr@  M;X
   court_hearrA  M<X   cousinrB  M=X   cranerC  M>X   crazyrD  M?X   crematerE  M@X
   cremationerF  MAX	   cresswellrG  MBX   cristalrH  MCX   crossingrI  MDX   croydonrJ  MEX
   cruiseboatrK  MFX   crusaderL  MGX   csirorM  MHX   cubanrN  MIX   culturerO  MJX   cuperrP  MKX   curtainrQ  MLX   curverR  MMX	   customaryrS  MNX   cyclewayrT  MOX   cyclistrU  MPX   dalbyrV  MQX   damnrW  MRX   dancerX  MSX   dangerrY  MTX	   dangerousrZ  MUX   darcyr[  MVX   darknessr\  MWX   darlingr]  MXX	   davenportr^  MYX   davyr_  MZX   dawesr`  M[X   dawkinra  M\X   dealerrb  M]X   deanrc  M^X   declarationrd  M_X
   defamationre  M`X   definerf  MaX	   deformityrg  MbX   defuserh  McX   defyri  MdX	   delightedrj  MeX   delugerk  MfX	   democracyrl  MgX	   dependentrm  MhX   depletern  MiX   depressro  MjX   derelictrp  MkX   designrq  MlX	   detectiverr  MmX   devonishrs  MnX   dialoguert  MoX   diamondru  MpX   dieselrv  MqX	   difficultrw  MrX   dilemmarx  MsX   dingory  MtX   dinnerrz  MuX	   directiver{  MvX   disabler|  MwX   disappointedr}  MxX   disappointingr~  MyX   disarmamentr  MzX	   discharger�  M{X   disciplinaryr�  M|X   discloser�  M}X   disconnectedr�  M~X   dismisser�  MX
   distributer�  M�X   distributorr�  M�X   diverr�  M�X   divingr�  M�X   dizzyr�  M�X   docklandr�  M�X   documentr�  M�X   doolanr�  M�X   doublyr�  M�X   downplayr�  M�X	   downshiftr�  M�X   downturnr�  M�X   downwardr�  M�X	   downwardsr�  M�X   draper�  M�X   drivingr�  M�X	   duckworthr�  M�X   dutyr�  M�X   eddysr�  M�X	   editorialr�  M�X   elderr�  M�X
   electronicr�  M�X   employr�  M�X   emptyr�  M�X   emulater�  M�X   endorser�  M�X   energyr�  M�X   engulfr�  M�X   enhancer�  M�X   enjoyr�  M�X
   enterpriser�  M�X   entertainmentr�  M�X   entrancer�  M�X   equalityr�  M�X	   eradicater�  M�X   errorr�  M�X
   evacuationr�  M�X	   eventuater�  M�X   evictr�  M�X   examinationr�  M�X   exceedr�  M�X	   excellentr�  M�X   existr�  M�X
   experiencer�  M�X   exploder�  M�X   extendedr�  M�X   extentr�  M�X   extinctr�  M�X
   extinctionr�  M�X   faceliftr�  M�X   fairfaxr�  M�X	   fareweller�  M�X   feastr�  M�X	   financingr�  M�X   firmr�  M�X
   fisichellar�  M�X   flamer�  M�X   flasherr�  M�X	   floodgater�  M�X   flushr�  M�X   fractionr�  M�X   freemanr�  M�X	   freighterr�  M�X   fridger�  M�X	   frustrater�  M�X   fudger�  M�X   fumer�  M�X   gadgetr�  M�X   gagr�  M�X   galleryr�  M�X   gazzar�  M�X   genuiner�  M�X   gingerr�  M�X   glitchr�  M�X
   governancer�  M�X   graduater�  M�X
   grandstandr�  M�X   graphicr�  M�X   grappler�  M�X   grassr�  M�X   graver�  M�X   grazingr�  M�X   grindr�  M�X   groomr�  M�X   grossr�  M�X   guitarr�  M�X   hammerr�  M�X   handedr�  M�X   happenr�  M�X   harassr�  M�X   hatchr�  M�X   hazardr�  M�X   headacher�  M�X	   headstoner�  M�X   helmetr�  M�X   heroer�  M�X   heroinr�  M�X   hijackr�  M�X   hiker�  M�X   hinderr�  M�X   homelandr�  M�X   homelessnessr�  M�X   hospitalisedr�  M�X   iconr�  M�X   imageryr�  M�X	   immigrantr�  M�X   immoralr�  M�X   inaugurationr�  M�X	   incorrectr�  M�X   independienter�  M�X   inflammatoryr�  M�X   influxr�  M�X   informationr�  M�X   initiater�  M�X
   initiativer�  M�X
   injunctionr�  M�X	   innocencer�  M�X   insider�  M�X   installationr�  M�X	   integrityr�  M�X	   intensifyr�  M�X	   intensityr�  M�X	   intentionr�  M�X   internalr   M�X
   internallyr  M�X	   intervener  M�X
   intimidater  M�X	   inventoryr  M�X
   invitationr  M X   involver  MX	   itinerantr  MX   joker  MX   jumperr	  MX   juniorr
  MX   jurorr  MX   kasperr  MX   keownr  MX
   kidnappingr  M	X   kingfishr  M
X   kniver  MX
   laboratoryr  MX   lakerr  MX   landminer  MX   languager  MX
   launderingr  MX   legislationr  MX
   legitimacyr  MX   leisurer  MX   lessenr  MX   liaisonr  MX   libertarianr  MX   lighterr  MX   limbor  MX   lingerr  MX   listenr  MX   loadingr   MX   lockr!  MX   lorientr"  MX   loverr#  MX   luckyr$  MX
   magistrater%  M X   magnetr&  M!X   magnificentr'  M"X   malaiser(  M#X   malariar)  M$X   manager*  M%X	   mandatoryr+  M&X   manhuntr,  M'X   manufacturer-  M(X   maroneyr.  M)X   maroochydorer/  M*X   marxistr0  M+X   massacrer1  M,X   massur2  M-X   mayr3  M.X   meatworkr4  M/X	   mediationr5  M0X   mercyr6  M1X
   microscoper7  M2X   migrater8  M3X	   migrationr9  M4X   militiar:  M5X   miner;  M6X   ministerialr<  M7X   mirrorr=  M8X   mistreatr>  M9X   modestr?  M:X	   molestingr@  M;X
   monitoringrA  M<X   moprB  M=X   morningrC  M>X   mortagerD  M?X   motloprE  M@X
   motorcrossrF  MAX   motorcyclistrG  MBX   mountainrH  MCX   moverrI  MDX   multinationalrJ  MEX   museeuwrK  MFX   muslimrL  MGX
   mysteriousrM  MHX   namibianrN  MIX
   neglectingrO  MJX	   negotiaterP  MKX   neighbourhoodrQ  MLX	   netballerrR  MMX   newbornrS  MNX	   northerlyrT  MOX   oasisrU  MPX   objectorrV  MQX   obscenerW  MRX   oceanrX  MSX   olympianrY  MTX   oneillrZ  MUX   onliner[  MVX   operater\  MWX   opinionr]  MXX   opportunityr^  MYX   oranger_  MZX   ordealr`  M[X   organra  M\X   organisationrb  M]X   orphanrc  M^X   outbackrd  M_X   outdoorsre  M`X   outlinerf  MaX   outrightrg  MbX   overambitiousrh  McX	   overbookeri  MdX   overlookrj  MeX	   overpowerrk  MfX   oysterrl  MgX
   pacesetterrm  MhX   paintingrn  MiX   pannero  MjX   paradornrp  MkX	   paralysedrq  MlX	   parameterrr  MmX   parishers  MnX   parkrt  MoX   parkingru  MpX   paroorv  MqX   passportrw  MrX   pastorrx  MsX   patriotry  MtX   patrolrz  MuX   pawnr{  MvX   payoutr|  MwX
   pedestrianr}  MxX   pegr~  MyX   pender  MzX	   penetrater�  M{X   pensionr�  M|X   petrol_pricer�  M}X
   philippiner�  M~X   phillipr�  MX   pileupr�  M�X   pillager�  M�X   pinpointr�  M�X   piper�  M�X   plainr�  M�X   plater�  M�X   playngr�  M�X
   playwrightr�  M�X
   plebisciter�  M�X   poacherr�  M�X   policewomanr�  M�X	   portfolior�  M�X   postalr�  M�X   postponementr�  M�X   pourr�  M�X   powellr�  M�X   preserver�  M�X   pressr�  M�X   pricingr�  M�X   priestr�  M�X   primer�  M�X	   principalr�  M�X   privacyr�  M�X   probablyr�  M�X   proceedr�  M�X
   processingr�  M�X   proclaimr�  M�X	   promisingr�  M�X   proner�  M�X   proteasr�  M�X   proudr�  M�X   providerr�  M�u(X   psychr�  M�X   pummelr�  M�X   pumpingr�  M�X   puncturer�  M�X   punterr�  M�X   purchaser�  M�X   putr�  M�X   puttingr�  M�X   quailr�  M�X
   queenslandr�  M�X   quicklyr�  M�X   quietr�  M�X   racingr�  M�X   rampantr�  M�X   ranger�  M�X   rangerr�  M�X   ratingr�  M�X	   readinessr�  M�X   realr�  M�X   rebater�  M�X   reboundr�  M�X	   receptionr�  M�X   reclaimr�  M�X   recommendationr�  M�X   recommendedr�  M�X   reconstructionr�  M�X   recreationalr�  M�X   recruitmentr�  M�X   redirectr�  M�X
   referendumr�  M�X   refineryr�  M�X	   refshauger�  M�X
   regulationr�  M�X	   reinstater�  M�X   reliancer�  M�X   relicr�  M�X
   relocationr�  M�X   remindr�  M�X   renaissancer�  M�X   renmarkr�  M�X
   renovationr�  M�X   rentalr�  M�X
   reportedlyr�  M�X   reporterr�  M�X   representationr�  M�X	   reprimandr�  M�X   rescuerr�  M�X   reserver�  M�X	   residencer�  M�X   respondr�  M�X   restedr�  M�X	   resurrectr�  M�X   resuscitationr�  M�X   reunificationr�  M�X   reuser�  M�X   rewardr�  M�X   ricochetr�  M�X
   ridiculousr�  M�X   riler�  M�X	   roadhouser�  M�X   robsonr�  M�X   rockyr�  M�X   romer�  M�X   roomr�  M�X   rotater�  M�X   rubbishr�  M�X   ruckerr�  M�X   ruinr�  M�X   sabrir�  M�X   sacredr�  M�X	   sacrificer�  M�X   salaryr�  M�X   scamr�  M�X   scammer�  M�X   scottishr�  M�X   selectr�  M�X   serenar�  M�X   sergeantr�  M�X   serialr�  M�X
   servicemanr�  M�X   sexualr�  M�X   shakyr�  M�X   shaper�  M�X   sharemarketr�  M�X   shatterr�  M�X   shedr�  M�X   shellr�  M�X   shelterr�  M�X   shiftr�  M�X   shoutr�  M�X   shrinkr�  M�X   significantr   M�X   silentr  M�X   sitterr  M�X   sixer  M�X   sixerr  M�X   sizer  M X	   skyrocketr  MX   slightlyr  MX   slugr  MX   smiler	  MX   solidr
  MX   soundr  MX	   sparinglyr  MX   spawningr  MX	   speculater  M	X   speedingr  M
X   spinalr  MX   spinnerr  MX   spitr  MX   sponsorr  MX   sponsorshipr  MX   springr  MX   sprintr  MX	   stanbroker  MX   stanwellr  MX   statr  MX   staunchr  MX   staver  MX   stickyr  MX   stifler  MX   stirr  MX	   stockpiler  MX   stormerr   MX
   strategistr!  MX   streamr"  MX   stretchr#  MX   strifer$  MX   stuffr%  M X	   subsidiser&  M!X   substandardr'  M"X   suburbr(  M#X
   successfulr)  M$X   suitabler*  M%X   sumr+  M&X   summerr,  M'X	   sunflowerr-  M(X   sunnierr.  M)X   superannuationr/  M*X	   superbiker0  M+X   surferr1  M,X   sustainr2  M-X   swansongr3  M.X   sweatr4  M/X   tamperr5  M0X   taskr6  M1X   tassiesr7  M2X   taster8  M3X   taxr9  M4X   teachingr:  M5X	   temporaryr;  M6X
   terminallyr<  M7X   thankfulr=  M8X   theatrer>  M9X	   thresholdr?  M:X   thunderr@  M;X   thwartrA  M<X   timidrB  M=X   tolerantrC  M>X   torchrD  M?X   torinorE  M@X	   tormentorrF  MAX   tottirG  MBX   toughenrH  MCX   towerrI  MDX   transparentrJ  MEX   traprK  MFX   trashrL  MGX   trendrM  MHX   trophierN  MIX   trouperO  MJX   tumourrP  MKX   turningrQ  MLX   umpirerR  MMX   unauthorisedrS  MNX   unavoidablerT  MOX   unawarerU  MPX   unconventionalrV  MQX	   underlinerW  MRX	   underminerX  MSX   unfencedrY  MTX	   universalrZ  MUX   universitier[  MVX   unsatisfactoryr\  MWX   unsolver]  MXX   upholdr^  MYX   uprisingr_  MZX   upstager`  M[X   urbanra  M\X   usualrb  M]X   vaguerc  M^X   valuerd  M_X   vampre  M`X	   vegetablerf  MaX   viewerrg  MbX   villierrh  McX	   violationri  MdX	   virtuallyrj  MeX   voicerk  MfX   volkerrl  MgX   warmingrm  MhX   warpathrn  MiX   wartimero  MjX   waywardrp  MkX   weakenrq  MlX   weaknessrr  MmX   wifers  MnX   willingrt  MoX   windfallru  MpX   windowrv  MqX   wineryrw  MrX   winterrx  MsX   witchry  MtX   withholdrz  MuX
   wollongongr{  MvX   wonderr|  MwX   workmanshipr}  MxX	   workplacer~  MyX   yieldr  MzX   youngestr�  M{X   abysmalr�  M|X   accommodationr�  M}X   accreditationr�  M~X   acquirer�  MX   additionr�  M�X	   advertiser�  M�X   afloatr�  M�X   alignr�  M�X	   allowancer�  M�X   alpolfor�  M�X   alreadyr�  M�X   amorusor�  M�X   amountr�  M�X   ankler�  M�X   anxietyr�  M�X   anzacr�  M�X   appallinglyr�  M�X
   appearancer�  M�X   appeaser�  M�X
   apprenticer�  M�X	   arrogancer�  M�X   attachr�  M�X
   attendancer�  M�X   attractr�  M�X   authorr�  M�X   avenuer�  M�X   backdownr�  M�X   baddeleyr�  M�X   bailr�  M�X	   ballisticr�  M�X   bankcardr�  M�X   barelyr�  M�X   barger�  M�X   barwonr�  M�X	   battalionr�  M�X   beaconr�  M�X	   behaviourr�  M�X   berthr�  M�X   billr�  M�X   binger�  M�X
   bipartisanr�  M�X   birthingr�  M�X   bloomr�  M�X   blowoutr�  M�X   blunderr�  M�X   boatier�  M�X   bondr�  M�X   boner�  M�X   bootr�  M�X   botanicr�  M�X   boundaryr�  M�X   bowlr�  M�X   boycottr�  M�X   branchr�  M�X	   brazilianr�  M�X   breakerr�  M�X   breastfeedingr�  M�X   breather�  M�X	   breathingr�  M�X   brickr�  M�X   britonr�  M�X   buggyr�  M�X   bunburyr�  M�X   bureaucracyr�  M�X	   burglarier�  M�X   bushlandr�  M�X   busyr�  M�X   cabinr�  M�X
   caboolturer�  M�X   calderr�  M�X   caltexr�  M�X   canior�  M�X   cannabir�  M�X   canningr�  M�X   canoer�  M�X   capellar�  M�X   capsicumr�  M�X   caravanr�  M�X   carryingr�  M�X
   cartoonistr�  M�X   caryardr�  M�X   cervicalr�  M�X   clarifier�  M�X   cliffr�  M�X   closedr�  M�X   cluer�  M�X
   collectionr�  M�X   columnr�  M�X   commandr�  M�X	   commodityr�  M�X   comparer�  M�X   competer�  M�X   concluder�  M�X
   confessionr�  M�X   confirmationr�  M�X   confuser�  M�X   conserver�  M�X   considerationr�  M�X   constitutionalr�  M�X
   constraintr�  M�X   contemplater�  M�X   contradictoryr�  M�X   controversyr�  M�X   conveniencer�  M�X   cooperativer�  M�X   copperr�  M�X   correctr�  M�X   corruptr�  M�X   costingr�  M�X   coughr�  M�X   countingr�  M�X   crabr�  M�X   craver�  M�X   crippledr�  M�X   crucifixionr�  M�X   crunchr�  M�X   cuffr�  M�X   curer�  M�X   cyclingr�  M�X   daisyr�  M�X   dancerr�  M�X   decader�  M�X   deciderr�  M�X   decreaser�  M�X   deedr�  M�X   deflectr�  M�X   demeritr�  M�X   demiser   M�X   demountabler  M�X   denialr  M�X   denmarkr  M�X   dentistr  M�X   deplorer  M X   deportationr  MX   derailr  MX
   derailmentr  MX
   deregulater	  MX   desperatelyr
  MX   detractr  MX
   difficultyr  MX   dirtyr  MX
   disabilityr  M	X	   disappearr  M
X   discardr  MX   disgracefulr  MX   distractr  MX   districtr  MX   ditchr  MX   dockingr  MX   doubtfulr  MX   downloadr  MX   downsizer  MX   dramar  MX   drillr  MX   drinkerr  MX   drinkingr  MX   droppingr  MX   drunkennessr  MX   easternr  MX   ecstasyr   MX   educater!  MX	   effectiver"  MX
   efficiencyr#  MX   ejectr$  MX
   electorater%  M X   electricr&  M!X   embarkr'  M"X
   embarrasser(  M#X   encircler)  M$X   enthroner*  M%X   entitler+  M&X   entrenchr,  M'X	   essentialr-  M(X   evaluater.  M)X   expirer/  M*X   explicitr0  M+X
   extinguishr1  M,X	   extortionr2  M-X   extraditionr3  M.X   failurer4  M/X   faithr5  M0X   falconerr6  M1X   fanningr7  M2X   fatallyr8  M3X   fellr9  M4X
   fellowshipr:  M5X   fingerr;  M6X   firearmr<  M7X   fitzroyr=  M8X   flanderr>  M9X   flarer?  M:X   flavorr@  M;X   floggingrA  M<X   foolishrB  M=X   footballrC  M>X   foretoldrD  M?X
   foundationrE  M@X   framerF  MAX   freakrG  MBX   fudgingrH  MCX   fuelrI  MDX   funnyrJ  MEX	   geriatricrK  MFX
   girlfriendrL  MGX   glarerM  MHX   gliderN  MIX   goldmanrO  MJX   goodrP  MKX   graftrQ  MLX	   guaranteerR  MMX   haemorrhagerS  MNX   handicaprT  MOX   hardwarerU  MPX   heatingrV  MQX   hesitantrW  MRX   highlyrX  MSX   higlightrY  MTX   hinklerrZ  MUX   hockeyr[  MVX   holdenr\  MWX
   honourabler]  MXX   horrifyr^  MYX   hotelierr_  MZX	   humiliater`  M[X   hussainra  M\X	   identifierb  M]X	   impendingrc  M^X   impersonaterd  M_X   implementationre  M`X	   implosionrf  MaX   impoundrg  MbX   inactionrh  McX	   inclusionri  MdX   incomingrj  MeX   inconclusiverk  MfX   independencerl  MgX   indictrm  MhX   infantrn  MiX   infectro  MjX   inflictrp  MkX	   injectionrq  MlX   inlandrr  MmX   insiderrs  MnX   inspectrt  MoX   insureru  MpX   intrv  MqX   intakerw  MrX   interconnectorrx  MsX	   interruptry  MtX   intersectionrz  MuX
   invaluabler{  MvX   involvedr|  MwX   irresponsibler}  MxX   jackr~  MyX   jackingr  MzX   jailedr�  M{X
   jeopardiser�  M|X   juventusr�  M}X   kiwir�  M~X   klimr�  MX   knockr�  M�X   ladenr�  M�X   landfillr�  M�X   laureater�  M�X   lawfulr�  M�X	   lawnmowerr�  M�X   leboucr�  M�X   lewdnessr�  M�X   libertadr�  M�X   limitedr�  M�X   locater�  M�X	   macarthurr�  M�X
   macfarlaner�  M�X	   machineryr�  M�X   mackayr�  M�X   mackerelr�  M�X   madridr�  M�X   magaziner�  M�X   magicr�  M�X   magicalr�  M�X   malpar�  M�X   mammalr�  M�X	   maralingar�  M�X   maritimer�  M�X	   marketingr�  M�X   marryr�  M�X   martynr�  M�X   masurr�  M�X   materr�  M�X   mccarthyr�  M�X   mcgradyr�  M�X   mcgraner�  M�X   mcguirer�  M�X   medicor�  M�X   mehrtenr�  M�X   mentorr�  M�X   meunierr�  M�X	   mgladbachr�  M�X   midwifer�  M�X   milanr�  M�X   millarr�  M�X   minardir�  M�X   misfirer�  M�X   moderater�  M�X   moleculer�  M�X   momentr�  M�X   monashr�  M�X   monsterr�  M�X
   montevideor�  M�X
   montgomeryr�  M�X   moochr�  M�X   mooneyr�  M�X   mortlockr�  M�X   moselyr�  M�X	   motocrossr�  M�X   motorr�  M�X   mournerr�  M�X   mulderr�  M�X   multiculturalr�  M�X   multipler�  M�X   mundiner�  M�X   muralr�  M�X
   murraylandr�  M�X   museumr�  M�X   mustardr�  M�X   muswellbrookr�  M�X   nacionalr�  M�X   nairnr�  M�X   nakedr�  M�X   nambourr�  M�X   nanter�  M�X   napler�  M�X   nattrassr�  M�X   naturer�  M�X
   naturopathr�  M�X	   necessaryr�  M�X   nedvedr�  M�X   nellyr�  M�X   nerver�  M�X   nervousr�  M�X   newlyr�  M�X
   newsagencyr�  M�X   nickelr�  M�X	   nightclubr�  M�X   nitschker�  M�X   noffker�  M�X
   nominationr�  M�X   noter�  M�X   noticer�  M�X   notifyr�  M�X   nuker�  M�X   nylexr�  M�X   obeidr�  M�X   observationr�  M�X   ofarrellr�  M�X	   offensiver�  M�X   oftenr�  M�X   ogradyr�  M�X   oilwellr�  M�X   oldfieldr�  M�X   olongar�  M�X   ominousr�  M�X   omissionr�  M�X   onesteelr�  M�X   ontarior�  M�X   organiser�  M�X	   organisedr�  M�X   orientationr�  M�X   originr�  M�X   osakar�  M�X	   osullivanr�  M�X   otherr�  M�X   ottenr�  M�X   otwayr�  M�X   outcomer�  M�X	   outnumberr�  M�X	   outspokenr�  M�X	   overspendr�  M�X   overworkr�  M�X	   ownershipr�  M�X	   pacemakerr�  M�X   paedophiliar�  M�X
   palaszczukr�  M�X   pamplingr   M�X   pantherr  M�X   parker  M�X	   parkinsonr  M�X   patiencer  M�X
   patriotismr  M X   patternr  MX   pauser  MX   penaliser  MX   penguinr	  MX	   peninsular
  MX   perkr  MX   permitr  MX   pettyr  MX   pharaohsr  M	X   pharmacyr  M
X   phialr  MX   photor  MX   photographerr  MX   pienaarr  MX   piercer  MX   pigeonr  MX   pigginr  MX   piperr  MX   piracyr  MX   pirer  MX   pirsar  MX   pitcairnr  MX   pittmanr  MX   pizzar  MX   playoffr  MX   pleasingr  MX   pocketr   MX   polishr!  MX   poochr"  MX   portraitr#  MX   portsear$  MX
   portsmouthr%  M X   potentr&  M!X   potentiallyr'  M"X   poultryr(  M#X   pozzator)  M$X
   pragmatismr*  M%X   prankr+  M&X   prattr,  M'X   preferr-  M(X	   prejudicer.  M)X   premeditater/  M*X   preselectionr0  M+X   primusr1  M,X	   processorr2  M-X	   profiteerr3  M.X   progr4  M/X	   promotionr5  M0X
   prospectorr6  M1X
   prostituter7  M2X   protear8  M3X	   publicityr9  M4X	   publisherr:  M5X   puckapunyalr;  M6X   pudder<  M7X   pumpr=  M8X   pursuitr>  M9X   pybusr?  M:X
   qantaslinkr@  M;X   queenslanderrA  M<X   questionablerB  M=X   questioningrC  M>X   racketrD  M?X   radarrE  M@X	   radclifferF  MAX	   radiationrG  MBX   railwayrH  MCX
   rainforestrI  MDX   rakerJ  MEX   ramsayrK  MFX   randomrL  MGX   rapperrM  MHX   ratificationrN  MIX   ratifyrO  MJX   rationaliserP  MKX	   ravanellirQ  MLX   ravensthorperR  MMX	   razorbackrS  MNX   reaffirmrT  MOX   receiverrU  MPX   recobarV  MQX   recyclerW  MRX	   redeveloprX  MSX   redundancierY  MTX   registrationrZ  MUX   regulater[  MVX	   regulatedr\  MWX   rehabr]  MXX   reignr^  MYX	   rejectionr_  MZX   rejuvenatedr`  M[X   relatera  M\X   relaxedrb  M]X   relegaterc  M^X
   relegationrd  M_X   remandre  M`X   remoterf  MaX	   renewablerg  MbX   reprieverh  McX   requirementri  MdX	   reservoirrj  MeX   respiterk  MfX
   restrainedrl  MgX   restrictiverm  MhX	   resurgentrn  MiX   reynoldro  MjX
   ricegrowerrp  MkX   riderrq  MlX   ridsdalerr  MmX   rigrs  MnX	   roadblockrt  MoX   roadsideru  MpX   robberyrv  MqX   robertrw  MrX   roddickrx  MsX   roederry  MtX   rosalindrz  MuX   roughingr{  MvX   routr|  MwX   roxbyr}  MxX   royaltyr~  MyX   ruffler  MzX   rushr�  M{X   sackingr�  M|X   saloonr�  M}X   sayyafr�  M~X	   schoolboyr�  MX
   schoolgirlr�  M�X	   schuttlerr�  M�X
   scientificr�  M�X   scornr�  M�X   scourger�  M�X   scrambler�  M�X   scrappedr�  M�X   scuffler�  M�X   seismicr�  M�X	   sensationr�  M�X   shipmentr�  M�X   shippingr�  M�X
   shoalhavenr�  M�X   shorer�  M�X	   shoreliner�  M�X   showier�  M�X   sideshowr�  M�X
   simplisticr�  M�X   singr�  M�X   singerr�  M�X	   situationr�  M�X	   skateparkr�  M�X   skittler�  M�X   slayr�  M�X   slightr�  M�X   snapperr�  M�X   sneakr�  M�X   snowyr�  M�X   snubr�  M�X   snuffr�  M�X   soberingr�  M�X   spikingr�  M�X   splurger�  M�X	   sportsbetr�  M�X   stallionr�  M�X   standardisationr�  M�X   standingr�  M�X   stanvacr�  M�X   steamr�  M�X	   steelworkr�  M�X   storer�  M�X   storyr�  M�X   strandedr�  M�X   strangerr�  M�X   stuartr�  M�X   stungr�  M�X   stuntr�  M�X   stuttler�  M�X   subduedr�  M�X	   substancer�  M�X   succumbr�  M�X   sudaneser�  M�X   suffererr�  M�X
   sunderlandr�  M�X	   supporterr�  M�X   surgicalr�  M�X	   surprisedr�  M�X   surveillancer�  M�X   switchr�  M�X   swordr�  M�X	   syndicater�  M�X   tallyr�  M�X   teachr�  M�X   tearr�  M�X   temporarilyr�  M�X   terrainr�  M�X   theoryr�  M�X   thinkerr�  M�X   throwerr�  M�X   thumpingr�  M�X   tiler�  M�X   timingr�  M�X   toiletr�  M�X	   tomahawksr�  M�X   toppler�  M�X   torpedor�  M�X   toutr�  M�X	   transformr�  M�X   trawlingr�  M�X	   triathlonr�  M�X   tshirtr�  M�X
   turnaroundr�  M�X   tussler�  M�X   twicer�  M�X   unacceptabler�  M�X
   undefeatedr�  M�X
   underwaterr�  M�X   unlawfulr�  M�X   unrulyr�  M�X   unsurprisedr�  M�X   unswayedr�  M�X   unwarrantedr�  M�X   uprootr�  M�X   user�  M�X   veerr�  M�X   verkerkr�  M�X   vigilr�  M�X   viker�  M�X   vitaminr�  M�X   voyager�  M�X   waltzr�  M�X   weakr�  M�X   webcastr�  M�X   websiter�  M�X   weedr�  M�X   weetwoodr�  M�X   wettestr�  M�X   whackr�  M�X	   wheatbeltr�  M�X   wherer�  M�X   willemr�  M�X   wingr�  M�X   workshopr�  M�X   worthr�  M�X   woundingr�  M�X   wrestler�  M�uX   id2tokenr�  }r�  X   cfsr�  }r�  (MKMKM�KM�KM�KM�KMK#M�KKMBK	M^KM;KMLKM�KM�KMVK
M KDK�KM�KM\K	M`KMRK	M!KM�K
M_KMEK:M�KM�KRMTKM]K3MKM�KM�KMbKKKBKMyK-M�KKTK-K�KM KMgKM�K	M�KMuK	M�KUMuKK	K4MyKK�K#M�KMKMEKM)KK�KM�K	M�KMKHM�MM~KKHKM�KMKM�K>MgKKKM�KMKM�KM[KMxK8MKKM�KM�K	M-KMKM�KMdKM-KK1KMIKMKMM�K}KKMcKMQKMkK
MjKM�KM�KMMKMUKKkK<M�KK�KMKMwKM<KVM�KKMUKEM�KM~KM_KM�KM1KK@KM�K	M�KM�KM�KM>KGM;KM�KM�KM�KIK
KM�K)K�KEMgKCK�KMFKMNKM�KDMKKMrKM@KMKMWKM�KM�KM�KMK
M�KM�KM�KM�KKFK	M#K=MbK MBKM�KMyKM�KMKKK)KMK9M�K/M�KM�K
M\KM{KMKMzKMKM�KK�K	K�KM�KM�KWM.KK�KKKKAKMwK2M�KMIK�MHK0M�K6M�KM5K�M.KMyK1MJK	MqKMfKMsK	M6KM�KM�KM%KMK0M=KM�K,M�KM�K
M�K+M�K	MKM1KM>K+M�KM�K M�KuM�KMKNMKM?KMyKIM�KM�KM�K"K,KK�K	M�KM�KMKK�K(M�K
M�KM)K;M"KM'KMdKMKM%KM#KM\K
M+KM�KM�KPM"KM�KM6KM@K	M�K%MGKM�K%MtKK�KMfKM�KM�KM3K3M1KM�K0M�KxM�KMiK�M�KMMKM�KM�KM�KM�KKKM�KM�KMIKM�KM.KM�KKDKM�KM
KK\K.M�KM�KM�KM�KM�KM�KM3K<MOKMQKMKK�KMUKMUK7MKM�KM�KM�KM�KM~KM�KM`KM)KM�K=M"KM�K'K�K M$KM�KM,KM:KM�KM=K/M�KMK)MZKMeKMeKK|K	K�KM�KM/KM8KM�K-MK'MXKM�KM�KMVKM�KMKM�KM�KM5KMKM�KMK"KLKKwKMvKMKMFKM�KM<K	M�K M�KM�K!M�K MdKMKBMKLMrKMqKM�KK�K'M[KM}KM|KM�KK.KKnKMuKK�KM4KKKK`KM\KM�KM�KMKK"KM�KM]KM�K8MWKMmKM�KM�KM�KMqKM@KM�KMKM�KM�KM	KM�KM1KM�KM�KMNKM`KMYKK!KM�K.M�KEM+KM�KM�K
KKMK
M.KMzKMVKMJK%KxKM�KMhKM�KMZKM�K	M�KM�KM�KM�K!M[K8M�KM�K	M�K;M0KMkKM`KM�K0MFKM0KM�KMKM.KM)KMKM�KM�KM�KjM�KM�KM@KM�KM�KKJKM�KMmKM~KM�KM�KM-KM�K
M�K-M�KM�KM KM�KM4KM�K
M�KM�KM�KM�KM�KM(KKMK
M�KMmKM�K
M�KMPK#M�KM*KMdK$MjK�M�KM�KM�KK{KK�K%MKMAKMvKM�KM�KM�KMK
M'KKKMfKMKM�KM�KM�KM�KMKMpKM�KM�KM�KM�KM�KMrKM�K!MwKM~KM�KMKK�KM�KK�KM�K3MOKM�KM6K	M>KM�KM�KMKMK$M
KM6KM�KKdKMfKMKM�KMEKM�KMDKM�KGMDKMFKMK MCK*M�KM�KK�KM7KK�KM�KM�KK+KM(KM�KM�KM�KM�KM�KM'KM~KMKMMK'KNKM�KMKMKM�KM�KM�KMKM�KM�KM�KMNKMiKM�KMkKK�KM#KM�K M�KK�KM�KGM2KMoKMzK&M"KM�KK�KMWKM�KM?KBM�K%M�K	MhKM%KMiKMnKM�KM�KM�KM,KMKMrKM�KGM{KM�K%K/KK�K*M�KMK	MKM�K/M�KM�KMOK*M�KM�K,K-K)M�K
M?KMhKMjKM�KM�KMBK	MNKM�KK�KOM�KK�KM�KMlKM K5MKM!KM5KMgKM�KM�KM�KMoKM�KM�KM�KM^KM>KM�KK�KMKMHKM�KM�KK>KM�KM�K1M�KM�K
MDKMSKM�KKgKMoKMK
M�KMKM�KM�KM�KM.KMWKMKM�KM�KKK+M�KMK K�KM�KM�KM1KM:KK�KM$K	MhKM�KMKM[KM�K	M�KBMtKM�KM KM�KM�KM�KM�KM�KM�K	M�KM�KMKM@KMKM�KM�K!MKKKM�KM#KM`KM8K"M+K5M�KMKM?KMqKM�KMlKM�KMKM�KM�K	M�KMKMtKM�K
M�KM�KMKM3K	M:KMKKM�KM&KM�KMrKK^KMBKM2KM�KK�KMKMtKM2KM�KMcK$M�KMjKM�KM�KMKM�KM�KM�KM_KM�KM'KM�KK�KMmKM�KM�KM�KM�KK:KMeKMvKM�KMOKKiKM�K#MeKK�KMOKM�KK KM�KM�KMyKM�KMKAM�KM�KMAKM=KM�K	M;K(KKMFKM|KM;KM�K:MJKK�KMKMKM�KKKMlKM�KMKM�KM�KM�KMZK	K�KM�KM�KM�KM�KM:KM�KM@KKKKKM�KM�KMKMSKM�K6M�KM�KMKM%KM�KMEK	M�K
M�K=MKM KM�KM�KM�K	M{KK�KM>KMQKM,KM	KMKMKMvKMLKKoKM�KM�K	KbKM�KM�KM�KM�KM#KMMKM�KM_KMlKMYKM�KM�KMzKM�KMtKM�KMMK
M}KM�K	M�KM�KMKKMPKMxKMKMK
M�KMyKMwK	M�KM
KM�KM�KM�KM%KM�KM�K%M2KM6KM�KMKM�K
M�KM�K"M�KK*KM:KMKM�KMYKKSKM�KK�KRM�KM�KKmKM�KM�KM�KM�KM�KSMxKMKM�KM�KM�KM<KoM�KM�KM?KK�KMfKK�KM�KM�KM�KK�KM�KM�KM,KM&KM9KMiKKKM�K.MwKM�KM�KM�KK&KMK!K�KM�KM�KM7KMKM�KM1KMZKM
K	M�K*M�KM�KM?KMqKMwKMKM�KMcKM�KK�KMKMK
M(KM�KM�KMKM�KM�KMaKK�KM�K	M�KM�KM�KM�KM�KMAKMmK6M'KMwK
MZK
M�KK�KMKMKM�KMKKKM�KMFKM�KMJKMGK&MWKMaKM=KM�KM�K
MpKM�KK�KKKK
MrKMKMGKMKM_KM9KM�KM+KMKMPKM�KM�K
M�KM�KM KMsKM�K(M(KMiKM�KMGKM�KM�KK#KM�KM�KM�KM�KM&KM KMjKMKM>KMEKM�KK7KM9KM�KMtKMKMcKK�Ku(K�K	M�KMK(MKM�K	M�K	M�KM�KKKMKM�KM�KMRKKhKM�KM�KK�KK8KMaKMHKMCKM�K	M8KM�KM�KM|KM�KM�KM�KMLKMGKMlKM�KM�KM�KK$KM�KM}KMKMKK�KM�KMKM\KMXKM�KM�KM�KM�KM�KMbKMKM$KK�K.M�KK�KMrKMdKMKM�KK�KM{KKKKRKMKM�KM�KM�KMCKM$KK�KKKMZKM%KMKM�KM�KK�KM�KM�K'MKMoKM�KKuKM�K	M0KK�KM0KM�KMZKM�K!M�KMXKM KM�KK;KK'KMKM�KMzKMKM�KK�KK�KM3KM^KM(KMBKM KMkKMKM�KMZKM�K'MKK�KM!KM�KMKM�KMKM�KM>KM�KM�KMnKM=KM7KK�KM-KMQKM}KK5KMKKKM\KM8KM�KM@KM�KMXKM�KKMKM�KMJKM�KM�KMuKM�K
M KMTKKKK�KM0KM�KM"KKK
M�KMeKMAK)MnKM�KM=K$MKMuKM�K	MKM�KK�KM�KM1KM�KM�KM4KMcKM�KM|KM�KM|KMKM�KM�KK�KM�KM�KM�KK�KM�KMKKKM�KM�KM�KK�KM�KM�KM�KMdKMcKM�KM�KM�KM�KM8KM)KKQKM
K
M�KMK
M]KM�K!MHKMKM�KM KMKM�KM�KM�KM�KMKM�K
K<KMQKK6KK�KM
KM�KM�KMKM�K(M�KMKM/KM�KMKM	KM�KM�KKfKM-KMKM�KM{KMXKM�KM�KM}KMRKM�KMxKM%KMK
M�K
KtKM�KM"KM�KM/KMKMvKMkKK�KM|KKeKM�KM�K	K_KM(KM�KM�KM<KM9KM�KM�KM�KK[KMNKM�KMKM�KM�KM)KM�K	M�KK�KM(K	M�KM�K	M�KM�KMGKK�KM�KMiKM�KMKM�KM/KMNKK=KM KM&KM�KM�KM�KM-KMHKM�KK�KMcKM�KKpKM+KM�K
KCKM�KK�KM�KMKM6KM�KMLKM�KMIKM�KMKM�KM4KM�KMIKM�KMUKM3KMaKMmKM�KMxKM�KM�KM�KM�KM*KM�KM	KMHKK�KM�KM�KM�KMDKMFKMPKMlKK�KM�KM�KMKM�KMVKMpKM�KM`KM�KK�KM�KMKM'KM=KM$KMhKK~KMKM]KMKMTKM;KM�KMMKM�KMeKM�KM@KM%KMaKM�KMJKM�KM�KK�KMzKMKM�KMbKMSK	M�KM�KM�KM�KM�KMKMVKMKMKMKKcK	M!KM�KK�KKKMsKM!KM�KM�KMpKM9K	MKM�KMKM.KMlKMKK�KMEKMeKK0KK�KM�KM�KM�KKYKMKM�KM{KM�KM�K	M�KM�KM�KM�KM�KK3KMEKMWKM
KM*KMKMDKM�KMKMUKMLKM�KM�KM}KMDKM�KMjKM�KM�KM�KKUKM�KM3KM�KK�KM�KM�KM�KM{KK�KMPKM�KMKM�KKrKM�KMYK
MKM�K
M�KMSKKVKMK	MuKK�KK�KM�KM�KM�KM�K	M�KM�KM�KM#KMKM�KM�KM�KM�KM�KMKM�KMKM!KK�KM&K
MKM$KMGKM9KK(KM�KM7KKIKM4KM�KMKM3KM�KM�KM�KMgKMzKM�KMKMgKMAKM�KM8KMfKK�KMKMKMYKM*KK9K
M�KMnKM�KM�KM�KM�KKGKM�KM�KMDKMxKM�KM�KM!KM�KMaKM�KMcKMmKM	KM�KM�KM�KMTKMNKMQKM�KM�KMKMWKM�K(K�KMKMsKM�KM+KM�KMKM*KMKMoKM�KM�KM�KM	KM2KM�KM[KM�KM�KM�KK�KM�KMtKM�KK�KKKK�KM�KMKMIKM�KM�KM�KM�KK�KM KMEKM7KM#KMQKM�KM�KM�KM�KK�KM�KM�KMvKMVKM|KM/KM�KKvK!K�KM�KMbKMKM4KMMKMqKK]KMbKM�KMMKM�KM�KMTKM5KM�KM�KMeKM;KM�KM�KM�KM�KM�KMKM�KM�KM�KMKMCKMKMXKMKM�KMKMRKM:KMKKMvKMvKMKM�KM\KM�K
MOKM�KM�K	M�KMKM�KKKM�KM~KM�KM�KMKMYKK�KM�KMXKM�KM'KMKMYKM^KM<K	MhKM�KM�KM�KM�KM�K
M�KMKM�K
M�KM�KMqKM�KMsKM�KM,KM�KM�KM�KM�KM�KM*KKjKM�KM�KMKM�KM�KM�KM5KMUKM�KMIKM�KM�KMaK
M6KM�KM�KM�KM�KMKM�KM�KM�KKyKM�KM�KM KM�KMKM�KMKMKM*KM�KM�KMKM�KM2KM�KMKM�KMCKM~KMKM�KK�KMhKM�KM[KM^KM�KM�KMpK	M^KMKM�KMKKK�KK�KM�KMkKM�KKzKM�KM8KM�KM�KMKMKM<KMKM7KMRKMOKM�KKKK�KM�KM�KM�KM�K	M3KMbKM1KM+KM�KMHKM�KM�KK�KMKMKMKM�KM�KM�KMkKMKMAKM2KM]KMhKK?KMbKMpKKEKMXKMKMjKM�KM�KM�KMuKMYK
M$KM�KM:KMnKM�KM�KM�KM�KM�KM�KM*KMKM�KMKM�KMLKM5KM�KMKM�KM�KM�KM5KMKM�KM�KM5KM�KM�KM(KM�KKsKMDKM�KM�KM)KM�KM�KK�KMmKMKM[KMxK
M�KKKM�KM�KM�KMLKM_KMK	M�KM<KMFKM&KM�KM�KMKKM�K	M�KMCKMKM�KMiKMKM�KMKM:KM�KMKKWKK�KKPKM�KM?KM�KM�KMHKM�KM!KM�KMBKM�KK�KK�KM&KM7KKaKM�KM>KMQKM�KM�KM�KMyKM{KM�KMCKM^KM|KM�KMoK MKM2KMdKMKM�KM'KM�KK�KMKMKM�KM�KM�KMVKM�KM)KMKM�KM\KMKM}K	K KM�KM�KM�KM?KMpKM4KMpKM�KM�KM�KM�KMKM0KM�KMkKM�KM�K	M�KMKM�KK�KMUKM-KM�KMKMKM�KMGKKlKMKM�K	M�KM�KM;KM�KM�KM�KM.KM�KMaKM0KK�KK�KM�KMoKK�KM�KMAKM,KM�KM�KMKM�Ku(MSKMtKM�KM;KM/KM�KM�KMoKMVKMjKM_KMTKKKM�KM/KM�KMsKMTKMLKMKM�KMJKM�KM�KMCKM�KK�KMKM7KM KM�KM�KK�KM�KMKM�KM�KMKM6KM�KM�KMKM�KM�KM�KMK
MKMPKM�KM`KM�KM�KM�KM�KM�KM�KKZKMBKM,KM�KMwKK%KK�KMRKM�KM8KM]KM�KM
KMSKM�KM�KM�KM�KM�KM�KM�KMnKMWKM�KM�KMKM9KMOKK�KMRKKOKM�KMuKMBKM�KM�KM+KM}KM�KM�KM�KM�KMqKM�KK�KM�KM`KM�KK}KM�KM�KKXKMSKM"KM/KM�KM$KMKMKM�KK�KM�KMKM-KMRKMPKM�KMfKK�KK�KMiKKKM4KM�KM#KK�KMfKMKM�KM�KM�KM�KM�KM�KM�K	K�KMnKM,KM�KM�KK�KM�KK�KM�KM�KMK	M�KK�KM0KM�KM�KM"KK�KMrKMgKMKM�KMKM]KMzKM�KMKM�KM_KK4KM�KMKM�KM�KM�KM�KM�KK�KM	KM=KM�KMnKM�KMgKM�K	M�KMsKM�KM�KKKMJKM�KM�KMPKMTKM�KMKK�KM&KM�KMlKM�KMKK�KM�KK�KM�KMNKM�KMSKK�KMIKM�KM�KMAKM�KM�KMKM�KMdKM�KM]KM�KMKMKM�KM<KM^KK2KM[KM�KK�KM	KM�KMKK�KM�KMxKMKM�KM�KKqKM�KM�KMKM9KM�KM�KM�KMsKM�KM�KM"	KMKMM
KM�KM�	KMF
KM�KM�	KMKMKM?KM8	KMGKM�K
M^KM�	KMKMeKM�KM�K!M�
KM�KM	KM�KM�KM�KM�KM	KM�KMKM'
KM�	KM�	KM�
KMM	KM|	KM�KM~	KMKKMK	MZKM�
KM�	KM�
KMhKM�	KM
KM�KM�	KM�
KMh
KM�KM�KM�	KM�KMg
KM�	KM�KM�	KM7KMKM	K
M�	KM3	KM�
KM�KMV
KM�KM�
KM�KM�	KM�KM�
KM�KM�	KM	KMVKM�KM�	KMNKM�KM(KM�
KM�KMX
KMKM�KM
KM1KM�	KMKM�	KM�	KM�	KMlKM�KM�KM�
KM�KM+
KM/KM
KMcKMUKMKMT	KMKM�KM�	KM6KM�KM�KM�KM�KM�	KMKM�KMsKM�KMY
KM-
KM�	KM�
KMJKM 
KM}KMW	KMHKM*	KM
KMKM�KM�KM�KMKM�	KM>KM�KM�KM�KMKM�KM>KMRKM�KM7
KMNKM
KM�	KM�KM4	KM�	KMm
KM;	KM�	KMhKM�
KMKM KM�KM�KM�	KM�
KMS
KMKM�KM`	KMd	KM@	KM�KM$KM�
KM9KM�
KM;KMKMLKMMKMKM�
KMBKM�	KM\KM�KM�
KM�
KM0	KM)KMKM�	KM KM�
KM�	KM
KM�KM�KMAKM�KMMKM�
KMzKM	KM�KMq	KMKM�
KMxKM`KM�KM<KM2	KM�KM�
KMi	KM�KM(
KMk	KM<	KM�KM;
KMO
KM�KM�KM�KM�KM%KM	KM�KMs
KM�KMKMKM1	KM�	KM5KM�KM]	KM
KM,KMpKM�	KM		KMvKM9	KM�KM
KMaKM�KM�KM
KM�KM KM�	KM�KM�
KM�	KM�KM�KM�
KM
KM�KM�KM�
KM�KM�
KM=
KMY	KMXKM�
KM�KMKM�
KMKM�	KMDKM�	KM:
KM�
KM]KM�KM�KM�
KM�KM�KM 	KMtKM�KM�KM$
KM5KM�
KM�KM�KM�
KMK	M�	KM	KMl
KMx
KM�KM#K	M�KM�
KMh	KM�
KM
KMUKMmKM�KM�	KMGKM`
KMKM|KM�KM�
KMKM�
KMl	KM�
KM�
KMn
KM
KM�KM�	KMQ	KM&KM�KM)
KM�	KM�
KM�KMX	KMz
KM�	KM�
KM8KM�	KM�	KM	KMKM3KM�KM8KM�KMf	KMCKMTKM^
KMb
KM`KMBKM�KM�KMKM�	KM�KM�KM�
KM�KM	KM�
KM�KM�	KMKMD
KM�KM�	KMyKM�KM�KM�KM	KM�KM�KM�KMsKM�	KM�KM�	KM�KMPKM�	KM�	KMzKM�
KM�KM:KM�KM�	KMqKM�KM:	KM�
KM�KM�	KMZ
KM�KM�
KM�KM�KM 	KM\
KM�
KM	KM	
KM&	KM�KM_KM/	KM	KM�KMKM�	KM�KMKMbKM�
KMJ
KMKM�	KM�	KM|
K
Mr
KM�KM�KM_KM�KM�
KMKMvKMm	KMlKMXKM
KM�KM�	KMKM�	KM�KM�KM7	KM�	KM�
KM_	KM�KM�
KM�KM�KM/KMU	KM<
KM�
KM�KM�
KM�KM�KM�KMKM�KMI
KM�KM	KM�KMRKM�KMv
KMWKM�	KM�
KMs	KMj
KM�	KM�KM�KMc	KM�KMx	KMKM6KM6	KM�
KMo
KMKM@KM
KM�KM	KM�KML	KM
KMD	KM0KM�	KML
KMYKM�KM&K
M�KME
KM4
KM�KM�	KM?
KM�
KM4KM�KM	KM�	KM	KM�KMq
KMw
KM)KM�
KM�
KM�KM�KMU
KMKMLKM�	KM�KM�KM�KM_
KM�KM�
KM�KMSKM�KM
KM�KM@KM�	KM,KM�KM�	KM2KM�KMg	KM�
KMR
KM�K
M�KM-KM�KM�KM�	KM�
KM!KM~KM;KM�KM�KM
KM�
KM	KMK	KM�KM�KMe
KMKM�
KM�
KM0KM	KM-	KM KM�
KMK
M�KMTKMKM�
KM	KM�KM�KM	KM�KM]KM,
KM3KM�KM�
KM�
KM
KM�
KMKM*KM[	KMA	KM�KM�
KM�	KMu	KM2KM�	KM�KMrKM�KM�
KM�KM	KMkKMKM�	KMa	KM�KM�
KM�KMy
KMKMwKMS	KM�
KM�KM�KM�KM�
KM�
KM�KM�KM!KM�KMn	KM
KM	KM�	KM
KM KM1KM�KM�KM�	KM�	KMnKM�
KM�K	MKM�KMnKM�KM�KMKMSKM�
KM�KM�	KMIKM#
KM7KM�KM�
KM6
KM�KM�KMP
KMoKM|KMIKM=KM[KM~
KM�KM�KM	KM�
KM�	KMKM�KMp
KM&
KMKM%	KMc
KM�KM�
KMKM*
KM�KMAKM�KMKM,	KMF	KM�KM	KM9KM�	KM�
KMKMG
KM�KM�KM-KM{	KMdKM�
KMwKM�	KMVKM�	KMj	KM�KM}	KM�
KM0
KM
KM
KMKMKM'KM\	KM�	KM
KM?	KMiKMp	KMxKM�	KMjKM�KM�KMWKM�KM�KM�
KM�
KMH	KM�KM{KM�	KM�
KM�
KM�KM�KM�	KMKM�	KMu
KM�	KM�KM�KM�KM�KM�	Ku(M�KM�KM�
KM�	KM.KM�KM�	KM"
KM]
KM�KM�KMFKM�	KM�KM�
KM	KM#KM�KM�KM�KMy	KM�
KMN	KM�
KMKM�KM�	KMKKM�	KM�
KM�	KM�KM�
KM 
KM)	KM!	KM�KM�KMt
KM�KM�KMf
KMgKMQKM$	KM�	KMN
KM�
KM	KMb	KM/
KMKM�	KMG	KMB
KM�KM�KM�KM{
KM�
KM	KMfKMi
KM[
KM9
KM}
KM�
KMqKM�	KM�
KM�	KM�KM�	KM�KM�KM�
KM�KM�KMQKM
KM
KM�
KM�
KM?KM�KM�KM�KM�	KM�
KM�KMKM�
KM�KM�KM�KM�
KM=KMKM�
KMoKM@
KM�KM	KM�	KM�KM(	KM�KM�	KMKM�
KM�KM'	KM�	KMuKM�	KM�
KM�	KMKMR	KM%
KM�KMKM�KM^	KM�KM�KM�KM�
KM�	KMJ	KM�	KM4KM�	KM�
KMFKM
KMuKMeKMv	KM5	KMKM	KM�
KM�KM�	KM�
KM�
KMP	KM�KMKM�	KMH
KM	KM�KM.
KM
	KMd
KMKM�	KMrKM�KMYKM
KM3
KMHKM2
KMK
KMmKM�
KM�	KM�	KM	KMk
KMaKM\KMe	KM�	KM
KM�KM�	KMQ
KM�
KM�KM^KM�	KM�	KM�KM*KMKM�KMKM�KM}KMJKMiKM"KM+	KMI	KM�KM�	KM�	KM�	KM�	KMEKM�KMKMKM%KM�KM�KMDKM�KM�KMa
KM�KM�KM.KM�
KM�KM�KM�KM�
KM�KM<KMt	KMyKM�KM�KM�K
M�KM�KMA
KM�
KM8
KMOKM�KM�KM�KMgKM�
KMbKM�
KMC	KMKM�KMO	KM"KM�KM~KM:KM�KM�
KM1
KM�KMr	KM�KMKMOKM'KM�	KM�KMZ	KM[KMjKM�KM�	KM>	KM.	KM�
KM#	KM!
KM�
KM�KM
KM�
KMPKM�
KM
KMC
KM{KM�
KM$KM�
KM�	KM�KM�KM�KM�KM�	KMtKM�KM�
KM�
KM	KM=	KMkKM�KM�KMB	KMfKMV	KMKM
KM�KM�KMcKM�	KM�
KM�KM�	KM�KM5
KMKMT
KM(KM+KM�KMKMZKM�
KM�KM	KM

KMW
KM�KMz	KMdKMw	KM�KM�	KMCKM
KMo	KMEKM>
KM�	KM�KM�KM
KM�KME	KM�	KMpKM�	KM+KM�KM^KM`KM2KM@KMeKMKM�KMrKMqKM�KM�KMKMKM�KM�KM-KM�KM�KM�KMCKM\KM�KM�KMcKMKMaKM�KMKMZKM.KM�KMiKM�KM*KM�KM1KM�KM'KM�KMUKM	KM�KMKM�KM�KMCKMKKM)KM=KM?KMhKMKMPKM�KMkKM�K	M^KM|KMKM-KM�KM�KM�KM9KM�KM�KM}KM#KMKM&KMzKM�KMCKMaKM�KMUKM�KM�KM�KMeKMZKMoKM�KM�KM�KM�KM2KM�KM'KMKM�KM�KMKM�KMpKM�KMKM�KMJKM�KM5KM$KMKM�KM�KM�KM~KM�KMcKMIKMXKM�KMgKM]KM"KMQKMVKM4KM�KMNKM�KM_KMfKMKM�KM�KMjKM�KM^KMWKMrKMcKMKM�KMuKM�KMKMRKMwK
M�KM�KM�KM�KM[KM�KMoKM]KM�KM�KM'KM$KMRKM�KMLKMKM>KMBKM�KMLKM8KM*KMGKMKM�KM&KM^KMuKM�KMPKM4KM�KM&KM+KM�KM�KM�KM�KM�KM�KM
KM`KM�KM�KMzKM KM�KM'KMXKM�KM�KMOKMIKM�KM�KM�KM�KMYKMDKM7KMlKMTKM�KM�KMKM�KM,KM�KM@KMAKM�KMDKM(KM�KM�KM?KM4KM�KM�KM0KM!KMKM�KMdKMFKM�KM"KMKM�KM�KMgKMJKMVKM�KMKM�KM~KM�KMSKMJKM�KMKMKMKM�KMWKMGKM�KM!KM�KMTKM[KMKM�KM�KM�KM�KM�KM�KM�KMxKM@KMKM�KMKMoKM*KMKMmKM�KMKMNKMKM6KM/KM�KM�KMKM�KM�KM1KMKMKMfKM�KM�KMkKM�KM�KMnKM�KM%KM5KMKMKM�KM�KMGKM�KMKM�KM_KMYKMKMkKMhKM�KM�KM�KM8KMKMKM�KM�KMqKMsKMvKM*KMoKM�KM~KM�KM�KM�KMKM�KM-KM1KM�KM�KM KM KM0KM5KMKMOKM�KMmKM�KM/KM8KM�KM�KMiKMmKM[KMKM�KM�KM�KMEKM�KM�KM�KMKM�KM}KMxKMyKM�KM�KMeKM�KMlKM:KM�KM�KMKM�KMHKM�KM�KM�KM,KM6KM�KMfKMcKMKKM9KMKM�KMKM`KM�KMYKM�KM�KMKMyKM=KM KMFKMUKM�KMhKMKMKM�KM�KMwKMDKM KM�KMdKM�KM�KMSKM�KMKMOKM�KMEKM�KMKM�KMpKMKM$KM�KMaKMzKM1KM�KM�KMWKM<KM(KM/KM�KMSKMKM.KM�KM[KMxKM�KMMKMBKM�KM�KM�KMKMBKM@KM�KM�KM�KM�KM�KM�KM�KM�KM�KM7KMKM�KM�KM�KMKM6KM�KMKM�KMdKM3KMMKMiKMsKMKM�KM�KM�KM�KM0KM�KM�KM�KMPKMDKM�KMZKMKM�KMKM:KMpKM�KM�KM�KM
KMvKM%KM�KM&KMKMqKM�KM3KM�KMVKM`KM�KMKM�KM.KM�KMGKMKM.KM�KMKM�KMKM$KM�KMEKMKM KMKM�KMnKM�KM�KMLKM]KM�KM�KM)KMeKM�KM�KM�KM�KM�KM�KMKMKM�KM�KM	KMKM>KM�KMMKM�KM�KMKMbKM>KM=KM�KM�KMKMWKM�KMKMbKM�KMiKM�KM�KM�KMKMZKM3KM	KM�KM�KM�KM�KMKM�KMIKM#KMxKM�KM]KM?KM�KM�KMKM%KMKM>KM�KM�KM�KMKKM�KMbKM�KM;KMtKMXKM�KM3KM�KMFKM�KMKM�KMwKM�KM�KM�KMKKM�KM�KM�KM�KM�KMCKM�KM�KM7KM�KM�KM"KM_KM�KM�KMYKM�KM�KMHKM�KM�KM�KM�KMXKMsKMgKMTKM\KMNKMBKM�KM9KM�KM;KM�KM?KM�KM�KM�KMMKMnKMIKM�KM�KMtKM�KM�KMOKu(M+KM�KM!KM�KMNKMHKMgKM,KMtKM�KM�KM<KM�KM�KM�KM2KM�KM�KM+KM�KM�KMKM�KMKM,KMKM/KM�KMmKM�KM�KMlKM�KM0KMuKMjKMlKM�KM�KMzKM�KM�KM-KMhKMKMfKM KM4KM%KMKM�KM�KM;KM#KMQKMEKMTKM�KMKMuKM�KMAKM;KM|KM�KM�KM+KMjKM�KM}KM�KM�KM�KM7KM�KM�KM�KMRKMAKMKM5KM�KM�KM�KM�KM(KM�KM�KMKM�KM�KMvKMKM�KM!KMQKM{KM�KM�KMaKM\KM�KM�KM�KMKMpKMKM�KM�KM8KM<KMAKM�KM�KM�KMdKMKM�KM"KM�KMKM�KM=KM�KM�KMKM�KM�KM�KM6KM�KMHKM�KM�KM�KM�KMvKM�KM�KM�KMnKM�KM:KM�KM�KM�KMqKM�KM�KMSKM�KMKM<KMJKM#KMFKMkKMQKMKM�KM�KM�KMPKM�KM:KM�KM�KM{KMjKMKM(KM�KM�KM�KMLKM_KM�KMrKM�KM�KM)KM�KMVKMwKMsKM�KM�KMKMKM�KM�KM�KMrKM�KMbKM9KMKMyKMUKMKM�KMKM{KM|KM
KM�KMKM{KMRKM2KM�KMtKMyKM�KMKM�KM�KMKM)KM\KM�KM�KMSKMKM�KMrKM�KM�KM�KM�KM�KMfKMKM�KM|KM�KM�KMoKM�KM�KM�KM�KMxKMqKM�KM�KM�KMKM�KM7KMWKM�KM�KMKM�KMKM�KM9KM8KM�KM�KM�KM�KM�KM!KM3KM�KM�KM�KM~KM�KMPKM�KM�KM�KMRKMxKM6KMuKM�KM�KM[KM�KMlKM�KM4KM�KMwKM�KM�KM�KMKM�KM�KM�KM�KM�KM�KM�KMKMsKM�KM�KMhKM�KM�KM�KM�KM+KM�KM�KM�KM5KMeKM�KMNKMKKMiKM�KM�KM�KMyKM�KM�KM�KM�KM=KMKMDKMKMRKM�KM`KM�KM�KMQKMLKMKM�KM�KM.KMZKM�KM�KM�KM�KM�KMjKMPKM�KM�KM KM�KM�KMBKM�KM?KM�KM�KMKM�KM�KMmKMHKMaKM�KM�KM�KMKMBKM�KM(KMVKM�KMHKM�KM�KM�KM�KM�KM%KMKMKMzKM�KMKM�KM�KM�KM�KM�KM�KM�KM�KMTKM
KM�KMiKM�KM�KM�KM�KM^KMhKMKMKMKM�KMYKM�KM1KM KM2KM�KM�KM�KM�KM�KM�KM�KM�KM}KMKM�KM�KM�KMFKM�KM�KM�KMuKMKM�KMbKM�KM�KMUKM�KMkKM�KM�KMIKM�KM�KM
KMXKM�KM�KM�KM�KM%KM�KM�KM�KM<KM�KM�KM.KM\KMMKM�KM�KMKMKMmKMNKM�KMrKM�KMdKM�KM�KM3KM�KMUKMKM�KM"KM�KM�KM�KM�KM�KM�KM�KM�KM!KM�KM�KM�KM�KMFKMKM;KMAKM�KMnKM_KM�KM�KM�KM�KM:KM�KMVKM�KMKM�KM�KM0KM�KMQKMqKM�KMIKM�KM}KM�KM�KMJKM�KM�KMOKMSKM,KM�KM�KM�KMGKM�KMfKM�KM�KM�KMJKM�KM�KM�KMKM8KM�KM~KM#KM�KM�KM�KM�KM�KM KM�KMKMKMKMpKMKM�KM�KM�KM�KM�KM�KM4KMvKM'KM�KM�KMKMgKM�KM_KM�KMKM�KM�KM KMcKM�KMWKMsKM�KM�KM,KMKM<KMoKM>KM�KM�KMcKMgKM�KM�KM`KM$KM�KMyKM)KMKM~KMKMvKMZKM�KM�KM6KM>KM�KMKM�KM�KM�KM�KM�KM"KM�KM(KM�KM�KM�KM�KM�KMTKM�KM�KM�KM�KM�KMLKM	KMKM�KM�KMXKM�KM*KM�KM�KM�KM}KM�KM�KM�KM�KM�KMKM�KM�KM�KMKM�KM�KM^KM'KM5KM�KM|KM�KM�KMYKM&KM[KMEKM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KMzKMKMtKM�KM�KM�KMdKM]KMnKM�KM?KM{KM�KM2KM�KM�KMKMKM�KMKM�KM�KM�KM�KMKKM�KMGKM\KM�KM|KM�KM�KMKMKM�KMDKM)KM�KM�KM�KM�KM�KM�KMKM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM/KM�KMKMCKM�KM1KM�KMOKM�KMKM�KM�KMKM�KMeKMKM&KM�KM=KM�KM�KM�KMEKM�KM�KM�KM	KM�KM:KM�KM@KM�KM�KM�KM�KM�KMKM�KMKM]KM�KM-KM7KM�KM�KM�KM�KM�KM�KM#KM�KM�KM�KM�KM�KM�KM�KM@KM�KM*KM�KM�KM�KM�KM�KMjKM;KM�KM�KMKMKM�KMKMCKM�KM�KM�KM0KMlKM�KMKM-KM�KM/KMkKM�KMKM�KM�KM�KMKMaKM$KM9KM�KM+KMKMKMwKM�KM�KM�KM�KM�KM�KM�KM�KMtKM�KMAKMbKM�KM�KM�KMKM�KM�KM{KM�KMpKMMKuX   dfsr�  }r�  (MKMKM�KM�KM�KM�KMKM�KMBKM^KM;KMLKM�KM�KMVKM KK�KM�KM\KM`KMRKM!KM�KM_KMEKM�KM�KMTKM]KMKM�KM�KMbKKBKMyKM�KKTKK�KM KMgKM�KM�KMuKM�KMuKK	KMyKK�KM�KMKMEKM)KK�KM�KM�KMKM�KM~KKHKM�KMKM�KMgKKKM�KMKM�KM[KMxKMKKM�KM�KM-KMKM�KMdKM-KK1KMIKMKM�KKKMcKMQKMkKMjKM�KM�KMMKMUKKkKM�KK�KMKMwKM<KM�KMUKM�KM~KM_KM�KM1KK@KM�KM�KM�KM�KM>KM;KM�KM�KM�KK
KM�KK�KMgKK�KMFKMNKM�KMKKMrKM@KMKMWKM�KM�KM�KMKM�KM�KM�KM�KKFKM#KMbKMBKM�KMyKM�KMKKK)KMKM�KM�KM�KM\KM{KMKMzKMKM�KK�KK�KM�KM�KM.KK�KKKKAKMwKM�KMIKMHKM�KM�KM5KM.KMyKMJKMqKMfKMsKM6KM�KM�KM%KMKM=KM�KM�KM�KM�KM�KMKM1KM>KM�KM�KM�KM�KMKMKM?KMyKM�KM�KM�KK,KK�KM�KM�KMKK�KM�KM�KM)KM"KM'KMdKMKM%KM#KM\KM+KM�KM�KM"KM�KM6KM@KM�KMGKM�KMtKK�KMfKM�KM�KM3KM1KM�KM�KM�KMiKM�KMMKM�KM�KM�KM�KKKM�KM�KMIKM�KM.KM�KKDKM�KM
KK\KM�KM�KM�KM�KM�KM�KM3KMOKMQKMKK�KMUKMUKMKM�KM�KM�KM�KM~KM�KM`KM)KM�KM"KM�KK�KM$KM�KM,KM:KM�KM=KM�KMKMZKMeKMeKK|KK�KM�KM/KM8KM�KMKMXKM�KM�KMVKM�KMKM�KM�KM5KMKM�KMKKLKKwKMvKMKMFKM�KM<KM�KM�KM�KM�KMdKMKMKMrKMqKM�KK�KM[KM}KM|KM�KK.KKnKMuKK�KM4KKKK`KM\KM�KM�KMKK"KM�KM]KM�KMWKMmKM�KM�KM�KMqKM@KM�KMKM�KM�KM	KM�KM1KM�KM�KMNKM`KMYKK!KM�KM�KM+KM�KM�KKKMKM.KMzKMVKMJKKxKM�KMhKM�KMZKM�KM�KM�KM�KM�KM[KM�KM�KM�KM0KMkKM`KM�KMFKM0KM�KMKM.KM)KMKM�KM�KM�KM�KM�KM@KM�KM�KKJKM�KMmKM~KM�KM�KM-KM�KM�KM�KM�KM KM�KM4KM�KM�KM�KM�KM�KM�KM(KMKM�KMmKM�KM�KMPKM�KM*KMdKMjKM�KM�KM�KK{KK�KMKMAKMvKM�KM�KM�KMKM'KKKMfKMKM�KM�KM�KM�KMKMpKM�KM�KM�KM�KM�KMrKM�KMwKM~KM�KMKK�KM�KK�KM�KMOKM�KM6KM>KM�KM�KMKMKM
KM6KM�KKdKMfKMKM�KMEKM�KMDKM�KMDKMFKMKMCKM�KM�KK�KM7KK�KM�KM�KK+KM(KM�KM�KM�KM�KM�KM'KM~KMKMMKKNKM�KMKMKM�KM�KM�KMKM�KM�KM�KMNKMiKM�KMkKK�KM#KM�KM�KK�KM�KM2KMoKMzKM"KM�KK�KMWKM�KM?KM�KM�KMhKM%KMiKMnKM�KM�KM�KM,KMKMrKM�KM{KM�KK/KK�KM�KMKMKM�KM�KM�KMOKM�KM�KK-KM�KM?KMhKMjKM�KM�KMBKMNKM�KK�KM�KK�KM�KMlKM KMKM!KM5KMgKM�KM�KM�KMoKM�KM�KM�KM^KM>KM�KK�KMKMHKM�KM�KK>KM�KM�KM�KM�KMDKMSKM�KKgKMoKMKM�KMKM�KM�KM�KM.KMWKMKM�KM�KKKM�KMKK�KM�KM�KM1KM:KK�KM$KMhKM�KMKM[KM�KM�KMtKM�KM KM�KM�KM�KM�KM�KM�KM�KM�KMKM@KMKM�KM�KMKKKM�KM#KM`KM8KM+KM�KMKM?KMqKM�KMlKM�KMKM�KM�KM�KMKMtKM�KM�KM�KMKM3KM:KMKKM�KM&KM�KMrKK^KMBKM2KM�KK�KMKMtKM2KM�KMcKM�KMjKM�KM�KMKM�KM�KM�KM_KM�KM'KM�KK�KMmKM�KM�KM�KM�KK:KMeKMvKM�KMOKKiKM�KMeKK�KMOKM�KK KM�KM�KMyKM�KMKM�KM�KMAKM=KM�KM;KKKMFKM|KM;KM�KMJKK�KMKMKM�KKKMlKM�KMKM�KM�KM�KMZKK�KM�KM�KM�KM�KM:KM�KM@KKKKKM�KM�KMKMSKM�KM�KM�KMKM%KM�KMEKM�KM�KMKM KM�KM�KM�KM{KK�KM>KMQKM,KM	KMKMKMvKMLKKoKM�KM�KKbKM�KM�KM�KM�KM#KMMKM�KM_KMlKMYKM�KM�KMzKM�KMtKM�KMMKM}KM�KM�KM�KMKKMPKMxKMKMKM�KMyKMwKM�KM
KM�KM�KM�KM%KM�KM�KM2KM6KM�KMKM�KM�KM�KM�KK*KM:KMKM�KMYKKSKM�KK�KM�KM�KKmKM�KM�KM�KM�KM�KMxKMKM�KM�KM�KM<KM�KM�KM?KK�KMfKK�KM�KM�KM�KK�KM�KM�KM,KM&KM9KMiKKKM�KMwKM�KM�KM�KK&KMKK�KM�KM�KM7KMKM�KM1KMZKM
KM�KM�KM�KM?KMqKMwKMKM�KMcKM�KK�KMKMKM(KM�KM�KMKM�KM�KMaKK�KM�KM�KM�KM�KM�KM�KMAKMmKM'KMwKMZKM�KK�KMKMKM�KMKKKM�KMFKM�KMJKMGKMWKMaKM=KM�KM�KMpKM�KK�KKKKMrKMKMGKMKM_KM9KM�KM+KMKMPKM�KM�KM�KM�KM KMsKM�KM(KMiKM�KMGKM�KM�KK#KM�KM�KM�KM�KM&KM KMjKMKM>KMEKM�KK7KM9KM�KMtKMKMcKK�Ku(K�KM�KMKMKM�KM�KM�KM�KKKMKM�KM�KMRKKhKM�KM�KK�KK8KMaKMHKMCKM�KM8KM�KM�KM|KM�KM�KM�KMLKMGKMlKM�KM�KM�KK$KM�KM}KMKMKK�KM�KMKM\KMXKM�KM�KM�KM�KM�KMbKMKM$KK�KM�KK�KMrKMdKMKM�KK�KM{KKKKRKMKM�KM�KM�KMCKM$KK�KKKMZKM%KMKM�KM�KK�KM�KM�KMKMoKM�KKuKM�KM0KK�KM0KM�KMZKM�KM�KMXKM KM�KK;KK'KMKM�KMzKMKM�KK�KK�KM3KM^KM(KMBKM KMkKMKM�KMZKM�KMKK�KM!KM�KMKM�KMKM�KM>KM�KM�KMnKM=KM7KK�KM-KMQKM}KK5KMKKKM\KM8KM�KM@KM�KMXKM�KKMKM�KMJKM�KM�KMuKM�KM KMTKKKK�KM0KM�KM"KKKM�KMeKMAKMnKM�KM=KMKMuKM�KMKM�KK�KM�KM1KM�KM�KM4KMcKM�KM|KM�KM|KMKM�KM�KK�KM�KM�KM�KK�KM�KMKKKM�KM�KM�KK�KM�KM�KM�KMdKMcKM�KM�KM�KM�KM8KM)KKQKM
KM�KMKM]KM�KMHKMKM�KM KMKM�KM�KM�KM�KMKM�KK<KMQKK6KK�KM
KM�KM�KMKM�KM�KMKM/KM�KMKM	KM�KM�KKfKM-KMKM�KM{KMXKM�KM�KM}KMRKM�KMxKM%KMKM�KKtKM�KM"KM�KM/KMKMvKMkKK�KM|KKeKM�KM�KK_KM(KM�KM�KM<KM9KM�KM�KM�KK[KMNKM�KMKM�KM�KM)KM�KM�KK�KM(KM�KM�KM�KM�KMGKK�KM�KMiKM�KMKM�KM/KMNKK=KM KM&KM�KM�KM�KM-KMHKM�KK�KMcKM�KKpKM+KM�KKCKM�KK�KM�KMKM6KM�KMLKM�KMIKM�KMKM�KM4KM�KMIKM�KMUKM3KMaKMmKM�KMxKM�KM�KM�KM�KM*KM�KM	KMHKK�KM�KM�KM�KMDKMFKMPKMlKK�KM�KM�KMKM�KMVKMpKM�KM`KM�KK�KM�KMKM'KM=KM$KMhKK~KMKM]KMKMTKM;KM�KMMKM�KMeKM�KM@KM%KMaKM�KMJKM�KM�KK�KMzKMKM�KMbKMSKM�KM�KM�KM�KM�KMKMVKMKMKMKKcKM!KM�KK�KKKMsKM!KM�KM�KMpKM9KMKM�KMKM.KMlKMKK�KMEKMeKK0KK�KM�KM�KM�KKYKMKM�KM{KM�KM�KM�KM�KM�KM�KM�KK3KMEKMWKM
KM*KMKMDKM�KMKMUKMLKM�KM�KM}KMDKM�KMjKM�KM�KM�KKUKM�KM3KM�KK�KM�KM�KM�KM{KK�KMPKM�KMKM�KKrKM�KMYKMKM�KM�KMSKKVKMKMuKK�KK�KM�KM�KM�KM�KM�KM�KM�KM#KMKM�KM�KM�KM�KM�KMKM�KMKM!KK�KM&KMKM$KMGKM9KK(KM�KM7KKIKM4KM�KMKM3KM�KM�KM�KMgKMzKM�KMKMgKMAKM�KM8KMfKK�KMKMKMYKM*KK9KM�KMnKM�KM�KM�KM�KKGKM�KM�KMDKMxKM�KM�KM!KM�KMaKM�KMcKMmKM	KM�KM�KM�KMTKMNKMQKM�KM�KMKMWKM�KK�KMKMsKM�KM+KM�KMKM*KMKMoKM�KM�KM�KM	KM2KM�KM[KM�KM�KM�KK�KM�KMtKM�KK�KKKK�KM�KMKMIKM�KM�KM�KM�KK�KM KMEKM7KM#KMQKM�KM�KM�KM�KK�KM�KM�KMvKMVKM|KM/KM�KKvKK�KM�KMbKMKM4KMMKMqKK]KMbKM�KMMKM�KM�KMTKM5KM�KM�KMeKM;KM�KM�KM�KM�KM�KMKM�KM�KM�KMKMCKMKMXKMKM�KMKMRKM:KMKKMvKMvKMKM�KM\KM�KMOKM�KM�KM�KMKM�KKKM�KM~KM�KM�KMKMYKK�KM�KMXKM�KM'KMKMYKM^KM<KMhKM�KM�KM�KM�KM�KM�KMKM�KM�KM�KMqKM�KMsKM�KM,KM�KM�KM�KM�KM�KM*KKjKM�KM�KMKM�KM�KM�KM5KMUKM�KMIKM�KM�KMaKM6KM�KM�KM�KM�KMKM�KM�KM�KKyKM�KM�KM KM�KMKM�KMKMKM*KM�KM�KMKM�KM2KM�KMKM�KMCKM~KMKM�KK�KMhKM�KM[KM^KM�KM�KMpKM^KMKM�KMKKK�KK�KM�KMkKM�KKzKM�KM8KM�KM�KMKMKM<KMKM7KMRKMOKM�KKKK�KM�KM�KM�KM�KM3KMbKM1KM+KM�KMHKM�KM�KK�KMKMKMKM�KM�KM�KMkKMKMAKM2KM]KMhKK?KMbKMpKKEKMXKMKMjKM�KM�KM�KMuKMYKM$KM�KM:KMnKM�KM�KM�KM�KM�KM�KM*KMKM�KMKM�KMLKM5KM�KMKM�KM�KM�KM5KMKM�KM�KM5KM�KM�KM(KM�KKsKMDKM�KM�KM)KM�KM�KK�KMmKMKM[KMxKM�KKKM�KM�KM�KMLKM_KMKM�KM<KMFKM&KM�KM�KMKKM�KM�KMCKMKM�KMiKMKM�KMKM:KM�KMKKWKK�KKPKM�KM?KM�KM�KMHKM�KM!KM�KMBKM�KK�KK�KM&KM7KKaKM�KM>KMQKM�KM�KM�KMyKM{KM�KMCKM^KM|KM�KMoKMKM2KMdKMKM�KM'KM�KK�KMKMKM�KM�KM�KMVKM�KM)KMKM�KM\KMKM}KK KM�KM�KM�KM?KMpKM4KMpKM�KM�KM�KM�KMKM0KM�KMkKM�KM�KM�KMKM�KK�KMUKM-KM�KMKMKM�KMGKKlKMKM�KM�KM�KM;KM�KM�KM�KM.KM�KMaKM0KK�KK�KM�KMoKK�KM�KMAKM,KM�KM�KMKM�Ku(MSKMtKM�KM;KM/KM�KM�KMoKMVKMjKM_KMTKKKM�KM/KM�KMsKMTKMLKMKM�KMJKM�KM�KMCKM�KK�KMKM7KM KM�KM�KK�KM�KMKM�KM�KMKM6KM�KM�KMKM�KM�KM�KMKMKMPKM�KM`KM�KM�KM�KM�KM�KM�KKZKMBKM,KM�KMwKK%KK�KMRKM�KM8KM]KM�KM
KMSKM�KM�KM�KM�KM�KM�KM�KMnKMWKM�KM�KMKM9KMOKK�KMRKKOKM�KMuKMBKM�KM�KM+KM}KM�KM�KM�KM�KMqKM�KK�KM�KM`KM�KK}KM�KM�KKXKMSKM"KM/KM�KM$KMKMKM�KK�KM�KMKM-KMRKMPKM�KMfKK�KK�KMiKKKM4KM�KM#KK�KMfKMKM�KM�KM�KM�KM�KM�KM�KK�KMnKM,KM�KM�KK�KM�KK�KM�KM�KMKM�KK�KM0KM�KM�KM"KK�KMrKMgKMKM�KMKM]KMzKM�KMKM�KM_KK4KM�KMKM�KM�KM�KM�KM�KK�KM	KM=KM�KMnKM�KMgKM�KM�KMsKM�KM�KKKMJKM�KM�KMPKMTKM�KMKK�KM&KM�KMlKM�KMKK�KM�KK�KM�KMNKM�KMSKK�KMIKM�KM�KMAKM�KM�KMKM�KMdKM�KM]KM�KMKMKM�KM<KM^KK2KM[KM�KK�KM	KM�KMKK�KM�KMxKMKM�KM�KKqKM�KM�KMKM9KM�KM�KM�KMsKM�KM�KM"	KMKMM
KM�KM�	KMF
KM�KM�	KMKMKM?KM8	KMGKM�KM^KM�	KMKMeKM�KM�KM�
KM�KM	KM�KM�KM�KM�KM	KM�KMKM'
KM�	KM�	KM�
KMM	KM|	KM�KM~	KMKKMKMZKM�
KM�	KM�
KMhKM�	KM
KM�KM�	KM�
KMh
KM�KM�KM�	KM�KMg
KM�	KM�KM�	KM7KMKM	KM�	KM3	KM�
KM�KMV
KM�KM�
KM�KM�	KM�KM�
KM�KM�	KM	KMVKM�KM�	KMNKM�KM(KM�
KM�KMX
KMKM�KM
KM1KM�	KMKM�	KM�	KM�	KMlKM�KM�KM�
KM�KM+
KM/KM
KMcKMUKMKMT	KMKM�KM�	KM6KM�KM�KM�KM�KM�	KMKM�KMsKM�KMY
KM-
KM�	KM�
KMJKM 
KM}KMW	KMHKM*	KM
KMKM�KM�KM�KMKM�	KM>KM�KM�KM�KMKM�KM>KMRKM�KM7
KMNKM
KM�	KM�KM4	KM�	KMm
KM;	KM�	KMhKM�
KMKM KM�KM�KM�	KM�
KMS
KMKM�KM`	KMd	KM@	KM�KM$KM�
KM9KM�
KM;KMKMLKMMKMKM�
KMBKM�	KM\KM�KM�
KM�
KM0	KM)KMKM�	KM KM�
KM�	KM
KM�KM�KMAKM�KMMKM�
KMzKM	KM�KMq	KMKM�
KMxKM`KM�KM<KM2	KM�KM�
KMi	KM�KM(
KMk	KM<	KM�KM;
KMO
KM�KM�KM�KM�KM%KM	KM�KMs
KM�KMKMKM1	KM�	KM5KM�KM]	KM
KM,KMpKM�	KM		KMvKM9	KM�KM
KMaKM�KM�KM
KM�KM KM�	KM�KM�
KM�	KM�KM�KM�
KM
KM�KM�KM�
KM�KM�
KM=
KMY	KMXKM�
KM�KMKM�
KMKM�	KMDKM�	KM:
KM�
KM]KM�KM�KM�
KM�KM�KM 	KMtKM�KM�KM$
KM5KM�
KM�KM�KM�
KMKM�	KM	KMl
KMx
KM�KM#KM�KM�
KMh	KM�
KM
KMUKMmKM�KM�	KMGKM`
KMKM|KM�KM�
KMKM�
KMl	KM�
KM�
KMn
KM
KM�KM�	KMQ	KM&KM�KM)
KM�	KM�
KM�KMX	KMz
KM�	KM�
KM8KM�	KM�	KM	KMKM3KM�KM8KM�KMf	KMCKMTKM^
KMb
KM`KMBKM�KM�KMKM�	KM�KM�KM�
KM�KM	KM�
KM�KM�	KMKMD
KM�KM�	KMyKM�KM�KM�KM	KM�KM�KM�KMsKM�	KM�KM�	KM�KMPKM�	KM�	KMzKM�
KM�KM:KM�KM�	KMqKM�KM:	KM�
KM�KM�	KMZ
KM�KM�
KM�KM�KM 	KM\
KM�
KM	KM	
KM&	KM�KM_KM/	KM	KM�KMKM�	KM�KMKMbKM�
KMJ
KMKM�	KM�	KM|
KMr
KM�KM�KM_KM�KM�
KMKMvKMm	KMlKMXKM
KM�KM�	KMKM�	KM�KM�KM7	KM�	KM�
KM_	KM�KM�
KM�KM�KM/KMU	KM<
KM�
KM�KM�
KM�KM�KM�KMKM�KMI
KM�KM	KM�KMRKM�KMv
KMWKM�	KM�
KMs	KMj
KM�	KM�KM�KMc	KM�KMx	KMKM6KM6	KM�
KMo
KMKM@KM
KM�KM	KM�KML	KM
KMD	KM0KM�	KML
KMYKM�KM&KM�KME
KM4
KM�KM�	KM?
KM�
KM4KM�KM	KM�	KM	KM�KMq
KMw
KM)KM�
KM�
KM�KM�KMU
KMKMLKM�	KM�KM�KM�KM_
KM�KM�
KM�KMSKM�KM
KM�KM@KM�	KM,KM�KM�	KM2KM�KMg	KM�
KMR
KM�KM�KM-KM�KM�KM�	KM�
KM!KM~KM;KM�KM�KM
KM�
KM	KMK	KM�KM�KMe
KMKM�
KM�
KM0KM	KM-	KM KM�
KMKM�KMTKMKM�
KM	KM�KM�KM	KM�KM]KM,
KM3KM�KM�
KM�
KM
KM�
KMKM*KM[	KMA	KM�KM�
KM�	KMu	KM2KM�	KM�KMrKM�KM�
KM�KM	KMkKMKM�	KMa	KM�KM�
KM�KMy
KMKMwKMS	KM�
KM�KM�KM�KM�
KM�
KM�KM�KM!KM�KMn	KM
KM	KM�	KM
KM KM1KM�KM�KM�	KM�	KMnKM�
KM�KMKM�KMnKM�KM�KMKMSKM�
KM�KM�	KMIKM#
KM7KM�KM�
KM6
KM�KM�KMP
KMoKM|KMIKM=KM[KM~
KM�KM�KM	KM�
KM�	KMKM�KMp
KM&
KMKM%	KMc
KM�KM�
KMKM*
KM�KMAKM�KMKM,	KMF	KM�KM	KM9KM�	KM�
KMKMG
KM�KM�KM-KM{	KMdKM�
KMwKM�	KMVKM�	KMj	KM�KM}	KM�
KM0
KM
KM
KMKMKM'KM\	KM�	KM
KM?	KMiKMp	KMxKM�	KMjKM�KM�KMWKM�KM�KM�
KM�
KMH	KM�KM{KM�	KM�
KM�
KM�KM�KM�	KMKM�	KMu
KM�	KM�KM�KM�KM�KM�	Ku(M�KM�KM�
KM�	KM.KM�KM�	KM"
KM]
KM�KM�KMFKM�	KM�KM�
KM	KM#KM�KM�KM�KMy	KM�
KMN	KM�
KMKM�KM�	KMKKM�	KM�
KM�	KM�KM�
KM 
KM)	KM!	KM�KM�KMt
KM�KM�KMf
KMgKMQKM$	KM�	KMN
KM�
KM	KMb	KM/
KMKM�	KMG	KMB
KM�KM�KM�KM{
KM�
KM	KMfKMi
KM[
KM9
KM}
KM�
KMqKM�	KM�
KM�	KM�KM�	KM�KM�KM�
KM�KM�KMQKM
KM
KM�
KM�
KM?KM�KM�KM�KM�	KM�
KM�KMKM�
KM�KM�KM�KM�
KM=KMKM�
KMoKM@
KM�KM	KM�	KM�KM(	KM�KM�	KMKM�
KM�KM'	KM�	KMuKM�	KM�
KM�	KMKMR	KM%
KM�KMKM�KM^	KM�KM�KM�KM�
KM�	KMJ	KM�	KM4KM�	KM�
KMFKM
KMuKMeKMv	KM5	KMKM	KM�
KM�KM�	KM�
KM�
KMP	KM�KMKM�	KMH
KM	KM�KM.
KM
	KMd
KMKM�	KMrKM�KMYKM
KM3
KMHKM2
KMK
KMmKM�
KM�	KM�	KM	KMk
KMaKM\KMe	KM�	KM
KM�KM�	KMQ
KM�
KM�KM^KM�	KM�	KM�KM*KMKM�KMKM�KM}KMJKMiKM"KM+	KMI	KM�KM�	KM�	KM�	KM�	KMEKM�KMKMKM%KM�KM�KMDKM�KM�KMa
KM�KM�KM.KM�
KM�KM�KM�KM�
KM�KM<KMt	KMyKM�KM�KM�KM�KM�KMA
KM�
KM8
KMOKM�KM�KM�KMgKM�
KMbKM�
KMC	KMKM�KMO	KM"KM�KM~KM:KM�KM�
KM1
KM�KMr	KM�KMKMOKM'KM�	KM�KMZ	KM[KMjKM�KM�	KM>	KM.	KM�
KM#	KM!
KM�
KM�KM
KM�
KMPKM�
KM
KMC
KM{KM�
KM$KM�
KM�	KM�KM�KM�KM�KM�	KMtKM�KM�
KM�
KM	KM=	KMkKM�KM�KMB	KMfKMV	KMKM
KM�KM�KMcKM�	KM�
KM�KM�	KM�KM5
KMKMT
KM(KM+KM�KMKMZKM�
KM�KM	KM

KMW
KM�KMz	KMdKMw	KM�KM�	KMCKM
KMo	KMEKM>
KM�	KM�KM�KM
KM�KME	KM�	KMpKM�	KM+KM�KM^KM`KM2KM@KMeKMKM�KMrKMqKM�KM�KMKMKM�KM�KM-KM�KM�KM�KMCKM\KM�KM�KMcKMKMaKM�KMKMZKM.KM�KMiKM�KM*KM�KM1KM�KM'KM�KMUKM	KM�KMKM�KM�KMCKMKKM)KM=KM?KMhKMKMPKM�KMkKM�KM^KM|KMKM-KM�KM�KM�KM9KM�KM�KM}KM#KMKM&KMzKM�KMCKMaKM�KMUKM�KM�KM�KMeKMZKMoKM�KM�KM�KM�KM2KM�KM'KMKM�KM�KMKM�KMpKM�KMKM�KMJKM�KM5KM$KMKM�KM�KM�KM~KM�KMcKMIKMXKM�KMgKM]KM"KMQKMVKM4KM�KMNKM�KM_KMfKMKM�KM�KMjKM�KM^KMWKMrKMcKMKM�KMuKM�KMKMRKMwKM�KM�KM�KM�KM[KM�KMoKM]KM�KM�KM'KM$KMRKM�KMLKMKM>KMBKM�KMLKM8KM*KMGKMKM�KM&KM^KMuKM�KMPKM4KM�KM&KM+KM�KM�KM�KM�KM�KM�KM
KM`KM�KM�KMzKM KM�KM'KMXKM�KM�KMOKMIKM�KM�KM�KM�KMYKMDKM7KMlKMTKM�KM�KMKM�KM,KM�KM@KMAKM�KMDKM(KM�KM�KM?KM4KM�KM�KM0KM!KMKM�KMdKMFKM�KM"KMKM�KM�KMgKMJKMVKM�KMKM�KM~KM�KMSKMJKM�KMKMKMKM�KMWKMGKM�KM!KM�KMTKM[KMKM�KM�KM�KM�KM�KM�KM�KMxKM@KMKM�KMKMoKM*KMKMmKM�KMKMNKMKM6KM/KM�KM�KMKM�KM�KM1KMKMKMfKM�KM�KMkKM�KM�KMnKM�KM%KM5KMKMKM�KM�KMGKM�KMKM�KM_KMYKMKMkKMhKM�KM�KM�KM8KMKMKM�KM�KMqKMsKMvKM*KMoKM�KM~KM�KM�KM�KMKM�KM-KM1KM�KM�KM KM KM0KM5KMKMOKM�KMmKM�KM/KM8KM�KM�KMiKMmKM[KMKM�KM�KM�KMEKM�KM�KM�KMKM�KM}KMxKMyKM�KM�KMeKM�KMlKM:KM�KM�KMKM�KMHKM�KM�KM�KM,KM6KM�KMfKMcKMKKM9KMKM�KMKM`KM�KMYKM�KM�KMKMyKM=KM KMFKMUKM�KMhKMKMKM�KM�KMwKMDKM KM�KMdKM�KM�KMSKM�KMKMOKM�KMEKM�KMKM�KMpKMKM$KM�KMaKMzKM1KM�KM�KMWKM<KM(KM/KM�KMSKMKM.KM�KM[KMxKM�KMMKMBKM�KM�KM�KMKMBKM@KM�KM�KM�KM�KM�KM�KM�KM�KM�KM7KMKM�KM�KM�KMKM6KM�KMKM�KMdKM3KMMKMiKMsKMKM�KM�KM�KM�KM0KM�KM�KM�KMPKMDKM�KMZKMKM�KMKM:KMpKM�KM�KM�KM
KMvKM%KM�KM&KMKMqKM�KM3KM�KMVKM`KM�KMKM�KM.KM�KMGKMKM.KM�KMKM�KMKM$KM�KMEKMKM KMKM�KMnKM�KM�KMLKM]KM�KM�KM)KMeKM�KM�KM�KM�KM�KM�KMKMKM�KM�KM	KMKM>KM�KMMKM�KM�KMKMbKM>KM=KM�KM�KMKMWKM�KMKMbKM�KMiKM�KM�KM�KMKMZKM3KM	KM�KM�KM�KM�KMKM�KMIKM#KMxKM�KM]KM?KM�KM�KMKM%KMKM>KM�KM�KM�KMKKM�KMbKM�KM;KMtKMXKM�KM3KM�KMFKM�KMKM�KMwKM�KM�KM�KMKKM�KM�KM�KM�KM�KMCKM�KM�KM7KM�KM�KM"KM_KM�KM�KMYKM�KM�KMHKM�KM�KM�KM�KMXKMsKMgKMTKM\KMNKMBKM�KM9KM�KM;KM�KM?KM�KM�KM�KMMKMnKMIKM�KM�KMtKM�KM�KMOKu(M+KM�KM!KM�KMNKMHKMgKM,KMtKM�KM�KM<KM�KM�KM�KM2KM�KM�KM+KM�KM�KMKM�KMKM,KMKM/KM�KMmKM�KM�KMlKM�KM0KMuKMjKMlKM�KM�KMzKM�KM�KM-KMhKMKMfKM KM4KM%KMKM�KM�KM;KM#KMQKMEKMTKM�KMKMuKM�KMAKM;KM|KM�KM�KM+KMjKM�KM}KM�KM�KM�KM7KM�KM�KM�KMRKMAKMKM5KM�KM�KM�KM�KM(KM�KM�KMKM�KM�KMvKMKM�KM!KMQKM{KM�KM�KMaKM\KM�KM�KM�KMKMpKMKM�KM�KM8KM<KMAKM�KM�KM�KMdKMKM�KM"KM�KMKM�KM=KM�KM�KMKM�KM�KM�KM6KM�KMHKM�KM�KM�KM�KMvKM�KM�KM�KMnKM�KM:KM�KM�KM�KMqKM�KM�KMSKM�KMKM<KMJKM#KMFKMkKMQKMKM�KM�KM�KMPKM�KM:KM�KM�KM{KMjKMKM(KM�KM�KM�KMLKM_KM�KMrKM�KM�KM)KM�KMVKMwKMsKM�KM�KMKMKM�KM�KM�KMrKM�KMbKM9KMKMyKMUKMKM�KMKM{KM|KM
KM�KMKM{KMRKM2KM�KMtKMyKM�KMKM�KM�KMKM)KM\KM�KM�KMSKMKM�KMrKM�KM�KM�KM�KM�KMfKMKM�KM|KM�KM�KMoKM�KM�KM�KM�KMxKMqKM�KM�KM�KMKM�KM7KMWKM�KM�KMKM�KMKM�KM9KM8KM�KM�KM�KM�KM�KM!KM3KM�KM�KM�KM~KM�KMPKM�KM�KM�KMRKMxKM6KMuKM�KM�KM[KM�KMlKM�KM4KM�KMwKM�KM�KM�KMKM�KM�KM�KM�KM�KM�KM�KMKMsKM�KM�KMhKM�KM�KM�KM�KM+KM�KM�KM�KM5KMeKM�KMNKMKKMiKM�KM�KM�KMyKM�KM�KM�KM�KM=KMKMDKMKMRKM�KM`KM�KM�KMQKMLKMKM�KM�KM.KMZKM�KM�KM�KM�KM�KMjKMPKM�KM�KM KM�KM�KMBKM�KM?KM�KM�KMKM�KM�KMmKMHKMaKM�KM�KM�KMKMBKM�KM(KMVKM�KMHKM�KM�KM�KM�KM�KM%KMKMKMzKM�KMKM�KM�KM�KM�KM�KM�KM�KM�KMTKM
KM�KMiKM�KM�KM�KM�KM^KMhKMKMKMKM�KMYKM�KM1KM KM2KM�KM�KM�KM�KM�KM�KM�KM�KM}KMKM�KM�KM�KMFKM�KM�KM�KMuKMKM�KMbKM�KM�KMUKM�KMkKM�KM�KMIKM�KM�KM
KMXKM�KM�KM�KM�KM%KM�KM�KM�KM<KM�KM�KM.KM\KMMKM�KM�KMKMKMmKMNKM�KMrKM�KMdKM�KM�KM3KM�KMUKMKM�KM"KM�KM�KM�KM�KM�KM�KM�KM�KM!KM�KM�KM�KM�KMFKMKM;KMAKM�KMnKM_KM�KM�KM�KM�KM:KM�KMVKM�KMKM�KM�KM0KM�KMQKMqKM�KMIKM�KM}KM�KM�KMJKM�KM�KMOKMSKM,KM�KM�KM�KMGKM�KMfKM�KM�KM�KMJKM�KM�KM�KMKM8KM�KM~KM#KM�KM�KM�KM�KM�KM KM�KMKMKMKMpKMKM�KM�KM�KM�KM�KM�KM4KMvKM'KM�KM�KMKMgKM�KM_KM�KMKM�KM�KM KMcKM�KMWKMsKM�KM�KM,KMKM<KMoKM>KM�KM�KMcKMgKM�KM�KM`KM$KM�KMyKM)KMKM~KMKMvKMZKM�KM�KM6KM>KM�KMKM�KM�KM�KM�KM�KM"KM�KM(KM�KM�KM�KM�KM�KMTKM�KM�KM�KM�KM�KMLKM	KMKM�KM�KMXKM�KM*KM�KM�KM�KM}KM�KM�KM�KM�KM�KMKM�KM�KM�KMKM�KM�KM^KM'KM5KM�KM|KM�KM�KMYKM&KM[KMEKM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KMzKMKMtKM�KM�KM�KMdKM]KMnKM�KM?KM{KM�KM2KM�KM�KMKMKM�KMKM�KM�KM�KM�KMKKM�KMGKM\KM�KM|KM�KM�KMKMKM�KMDKM)KM�KM�KM�KM�KM�KM�KMKM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM�KM/KM�KMKMCKM�KM1KM�KMOKM�KMKM�KM�KMKM�KMeKMKM&KM�KM=KM�KM�KM�KMEKM�KM�KM�KM	KM�KM:KM�KM@KM�KM�KM�KM�KM�KMKM�KMKM]KM�KM-KM7KM�KM�KM�KM�KM�KM�KM#KM�KM�KM�KM�KM�KM�KM�KM@KM�KM*KM�KM�KM�KM�KM�KMjKM;KM�KM�KMKMKM�KMKMCKM�KM�KM�KM0KMlKM�KMKM-KM�KM/KMkKM�KMKM�KM�KM�KMKMaKM$KM9KM�KM+KMKMKMwKM�KM�KM�KM�KM�KM�KM�KM�KMtKM�KMAKMbKM�KM�KM�KMKM�KM�KM{KM�KMpKMMKuX   num_docsr�  KX   num_posr   MGdX   num_nnzr  M�#X   __numpysr  ]r  X   __scipysr  ]r  X
   __ignoredsr  ]r  X   __recursive_saveloadsr  ]r	  ub.